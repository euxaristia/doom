module core

pub fn f_responder(ev &Event) bool {
	_ = ev
	return false
}

pub fn f_ticker() {}
pub fn f_drawer() {}
pub fn f_start_finale() {}
