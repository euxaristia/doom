module core

pub fn deh_doom_init() {}
