@[has_globals]
module core

__global deh_bex_strings_loaded = false

pub fn deh_bexstr_init() {
	deh_bex_strings_loaded = false
}
