@[translated]
module main

// Setup textscreen key input module: placeholder manual port.
