module core

pub fn deh_sound_init() {}
