@[translated]
module main

// V dehacked init shim: placeholder manual port.
