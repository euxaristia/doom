module core

pub fn p_plats_do_plat_stub(line &Line, plattype int, amount int) int {
	_ = line
	_ = plattype
	_ = amount
	return 0
}

pub fn p_plats_activate_in_stasis_stub(tag int) {
	_ = tag
}
