@[translated]
module main

// Textscreen input box widget: placeholder manual port.
