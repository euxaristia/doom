@[translated]
module main

// Textscreen conditional widget: placeholder manual port.
