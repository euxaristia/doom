module core

pub fn stat_copy(stats &WbStartStruct) {
	_ = stats
}

pub fn stat_dump() {}
