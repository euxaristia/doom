@[has_globals]
module core

pub const skyflatname = 'F_SKY1'
pub const angletoskyshift = 22

__global skytexture = 0
__global skytexturemid = 0

pub fn r_init_sky_map() {}
