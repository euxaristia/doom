@[has_globals]
module core

__global gameaction = GameAction.nothing

pub fn d_process_events() {
}

pub fn d_page_ticker() {
}

pub fn d_page_drawer() {
}

pub fn d_advance_demo() {
}

pub fn d_do_advance_demo() {
}

pub fn d_start_title() {
}
