@[translated]
module main

// Loopback networking support: placeholder manual port.
