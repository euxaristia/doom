@[has_globals]
module core

__global deh_ammo_overrides = 0

pub fn deh_ammo_init() {
	deh_ammo_overrides = 0
}
