@[translated]
module main

// Textscreen GUI test example: placeholder manual port.
