@[translated]
module main

// SDL networking support: placeholder manual port.
