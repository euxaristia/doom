@[translated]
module main

// Textscreen desktop widget: placeholder manual port.
