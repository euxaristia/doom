@[translated]
module main

// Networking client: placeholder manual port.
