@[translated]
module main

// SDL sound backend: placeholder manual port.
