@[translated]
module main

// Textscreen label widget: placeholder manual port.
