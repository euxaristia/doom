@[translated]
module main

// Textscreen table widget: placeholder manual port.
