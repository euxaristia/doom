module core

pub const savegamename = 'doomsav'
pub const num_quitmessages = 8

pub const doom1_endmsg = [
	'please do not leave',
	'you are a hero',
	'try again soon',
	'doom awaits',
	'monsters miss you',
	'one more level',
	'keep fragging',
	'farewell marine',
]

pub const doom2_endmsg = [
	'doom2 says bye',
	'no rest for you',
	'hell stays open',
	'come back armed',
	'you know the way',
	'still not enough',
	'just one more',
	'goodbye marine',
]
