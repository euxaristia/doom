@[translated]
module main

// Textscreen checkbox widget: placeholder manual port.
