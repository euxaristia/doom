@[translated]
module main

// Textscreen window action widget: placeholder manual port.
