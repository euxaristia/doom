@[translated]
module main

// Textscreen I/O module: placeholder manual port.
