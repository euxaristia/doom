module core

// Minimal renderer state placeholders.
pub fn r_init_state() {}
