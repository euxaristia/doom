@[translated]
module main

// Textscreen window widget: placeholder manual port.
