@[translated]
module main

// OPL queue: placeholder manual port.
