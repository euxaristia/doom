module core

// Enemy AI is not ported yet; keep entrypoints present.
pub fn p_enemy_think(mobj &Mobj) {
	_ = mobj
}

pub fn p_spawn_brain_targets() {}
pub fn p_clear_brain_targets() {}
