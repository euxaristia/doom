module core

pub fn r_render_segs() {}

pub fn r_render_masked_seg_range(ds &DrawSeg, x1 int, x2 int) {
	_ = ds
	_ = x1
	_ = x2
}
