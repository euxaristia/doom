@[translated]
module main

// Textscreen radio button widget: placeholder manual port.
