module core

// Renderer umbrella header placeholder.
pub fn r_init_local() {}
