@[translated]
module main

// Setup textscreen joystick button input module: placeholder manual port.
