@[translated]
module main

// Setup joystick module: placeholder manual port.
