@[translated]
module main

// OPL core: placeholder manual port.
