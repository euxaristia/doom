module core

pub struct Pic {
pub mut:
	width  u8
	height u8
	data   u8
}
