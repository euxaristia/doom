@[translated]
module main

// Setup textscreen mouse input module: placeholder manual port.
