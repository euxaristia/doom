module core

pub fn p_switch_change_texture_stub(line &Line, use_again int) {
	_ = line
	_ = use_again
}

pub fn p_switch_use_special_line_stub(mobj &Mobj, line &Line, side int) bool {
	_ = mobj
	_ = line
	_ = side
	return false
}
