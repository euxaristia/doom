@[translated]
module main

// Textscreen SDL backend: placeholder manual port.
