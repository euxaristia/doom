module core

pub fn deh_bexstr_init() {}
