module core

pub fn ev_teleport(line &Line, side int, thing &Mobj) int {
	_ = line
	_ = side
	_ = thing
	return 0
}
