module core

pub fn deh_thing_init() {}
