@[translated]
module main

// Win32 opendir compatibility: placeholder manual port.
