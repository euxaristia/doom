module core

pub fn p_check_sight_stub(t1 &Mobj, t2 &Mobj) bool {
	return p_check_sight(t1, t2)
}
