@[translated]
module main

// POSIX WAD file backend: placeholder manual port.
