@[translated]
module main

// Win32 WAD file backend: placeholder manual port.
