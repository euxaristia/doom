@[translated]
module main

// Setup multiplayer module: placeholder manual port.
