module core

pub fn deh_cheat_init() {}
