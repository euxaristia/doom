@[translated]
module main

// Network server support: placeholder manual port.
