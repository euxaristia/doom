module core

pub enum WiStateEnum {
	no_state = -1
	stat_count
	show_next_loc
}

pub fn wi_ticker() {}
pub fn wi_drawer() {}
pub fn wi_start(wbstartstruct &WbStartStruct) { _ = wbstartstruct }
pub fn wi_end() {}
