@[translated]
module main

// Network query support: placeholder manual port.
