module core

pub fn ev_do_floor(line &Line, floortype int) int {
	_ = line
	_ = floortype
	return 0
}
