module core

pub fn deh_ammo_init() {}
