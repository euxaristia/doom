@[translated]
module main

fn C.W_Init()
fn C.W_AutoLoad()
fn C.W_LoadRemainingLumps()

fn w_init() { C.W_Init() }
fn w_auto_load() { C.W_AutoLoad() }
fn w_load_remaining_lumps() { C.W_LoadRemainingLumps() }
