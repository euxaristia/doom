module core

// Placeholder tables module used by renderer headers.
pub const fine_angles = 8192
pub const fine_mask = fine_angles - 1

pub const finesine = []Fixed{}
pub const finecosine = []Fixed{}
