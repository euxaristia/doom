@[has_globals]
module core

__global deh_doom_loaded = false

pub fn deh_doom_init() {
	deh_doom_loaded = false
}
