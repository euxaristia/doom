module core

pub fn deh_ptr_init() {}
