@[has_globals]
module core

__global deh_ptr_overrides = 0

pub fn deh_ptr_init() {
	deh_ptr_overrides = 0
}
