@[translated]
module main

// Textscreen widget core: placeholder manual port.
