@[translated]
module main

// Textscreen scrollpane widget: placeholder manual port.
