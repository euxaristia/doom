module tables

@[translated]

const slope_range = 4096

fn slope_div(num u32, den u32) u32 {
    if den < 512 {
        return slope_range
    } else {
        ans := (num << 3) / (den >> 8)
        if ans <= slope_range {
            return ans
        } else {
            return slope_range
        }
    }
}

const finetangent = [i32(
-170910304,-56965752,-34178904,-24413316,-18988036,-15535599,-13145455,-11392683,
    -10052327,-8994149,-8137527,-7429880,-6835455,-6329090,-5892567,-5512368,
    -5178251,-4882318,-4618375,-4381502,-4167737,-3973855,-3797206,-3635590,
    -3487165,-3350381,-3223918,-3106651,-2997613,-2895966,-2800983,-2712030,
    -2628549,-2550052,-2476104,-2406322,-2340362,-2277919,-2218719,-2162516,
    -2109087,-2058233,-2009771,-1963536,-1919378,-1877161,-1836758,-1798063,
    -1760956,-1725348,-1691149,-1658278,-1626658,-1596220,-1566898,-1538632,
    -1511367,-1485049,-1459630,-1435065,-1411312,-1388330,-1366084,-1344537,
    -1323658,-1303416,-1283783,-1264730,-1246234,-1228269,-1210813,-1193846,
    -1177345,-1161294,-1145673,-1130465,-1115654,-1101225,-1087164,-1073455,
    -1060087,-1047046,-1034322,-1021901,-1009774,-997931,-986361,-975054,
    -964003,-953199,-942633,-932298,-922186,-912289,-902602,-893117,
    -883829,-874730,-865817,-857081,-848520,-840127,-831898,-823827,
    -815910,-808143,-800521,-793041,-785699,-778490,-771411,-764460,
    -757631,-750922,-744331,-737853,-731486,-725227,-719074,-713023,
    -707072,-701219,-695462,-689797,-684223,-678737,-673338,-668024,
    -662792,-657640,-652568,-647572,-642651,-637803,-633028,-628323,
    -623686,-619117,-614613,-610174,-605798,-601483,-597229,-593033,
    -588896,-584815,-580789,-576818,-572901,-569035,-565221,-561456,
    -557741,-554074,-550455,-546881,-543354,-539870,-536431,-533034,
    -529680,-526366,-523094,-519861,-516667,-513512,-510394,-507313,
    -504269,-501261,-498287,-495348,-492443,-489571,-486732,-483925,
    -481150,-478406,-475692,-473009,-470355,-467730,-465133,-462565,
    -460024,-457511,-455024,-452564,-450129,-447720,-445337,-442978,
    -440643,-438332,-436045,-433781,-431540,-429321,-427125,-424951,
    -422798,-420666,-418555,-416465,-414395,-412344,-410314,-408303,
    -406311,-404338,-402384,-400448,-398530,-396630,-394747,-392882,
    -391034,-389202,-387387,-385589,-383807,-382040,-380290,-378555,
    -376835,-375130,-373440,-371765,-370105,-368459,-366826,-365208,
    -363604,-362013,-360436,-358872,-357321,-355783,-354257,-352744,
    -351244,-349756,-348280,-346816,-345364,-343924,-342495,-341078,
    -339671,-338276,-336892,-335519,-334157,-332805,-331464,-330133,
    -328812,-327502,-326201,-324910,-323629,-322358,-321097,-319844,
    -318601,-317368,-316143,-314928,-313721,-312524,-311335,-310154,
    -308983,-307819,-306664,-305517,-304379,-303248,-302126,-301011,
    -299904,-298805,-297714,-296630,-295554,-294485,-293423,-292369,
    -291322,-290282,-289249,-288223,-287204,-286192,-285186,-284188,
    -283195,-282210,-281231,-280258,-279292,-278332,-277378,-276430,
    -275489,-274553,-273624,-272700,-271782,-270871,-269965,-269064,
    -268169,-267280,-266397,-265519,-264646,-263779,-262917,-262060,
    -261209,-260363,-259522,-258686,-257855,-257029,-256208,-255392,
    -254581,-253774,-252973,-252176,-251384,-250596,-249813,-249035,
    -248261,-247492,-246727,-245966,-245210,-244458,-243711,-242967,
    -242228,-241493,-240763,-240036,-239314,-238595,-237881,-237170,
    -236463,-235761,-235062,-234367,-233676,-232988,-232304,-231624,
    -230948,-230275,-229606,-228941,-228279,-227621,-226966,-226314,
    -225666,-225022,-224381,-223743,-223108,-222477,-221849,-221225,
    -220603,-219985,-219370,-218758,-218149,-217544,-216941,-216341,
    -215745,-215151,-214561,-213973,-213389,-212807,-212228,-211652,
    -211079,-210509,-209941,-209376,-208815,-208255,-207699,-207145,
    -206594,-206045,-205500,-204956,-204416,-203878,-203342,-202809,
    -202279,-201751,-201226,-200703,-200182,-199664,-199149,-198636,
    -198125,-197616,-197110,-196606,-196105,-195606,-195109,-194614,
    -194122,-193631,-193143,-192658,-192174,-191693,-191213,-190736,
    -190261,-189789,-189318,-188849,-188382,-187918,-187455,-186995,
    -186536,-186080,-185625,-185173,-184722,-184274,-183827,-183382,
    -182939,-182498,-182059,-181622,-181186,-180753,-180321,-179891,
    -179463,-179037,-178612,-178190,-177769,-177349,-176932,-176516,
    -176102,-175690,-175279,-174870,-174463,-174057,-173653,-173251,
    -172850,-172451,-172053,-171657,-171263,-170870,-170479,-170089,
    -169701,-169315,-168930,-168546,-168164,-167784,-167405,-167027,
    -166651,-166277,-165904,-165532,-165162,-164793,-164426,-164060,
    -163695,-163332,-162970,-162610,-162251,-161893,-161537,-161182,
    -160828,-160476,-160125,-159775,-159427,-159079,-158734,-158389,
    -158046,-157704,-157363,-157024,-156686,-156349,-156013,-155678,
    -155345,-155013,-154682,-154352,-154024,-153697,-153370,-153045,
    -152722,-152399,-152077,-151757,-151438,-151120,-150803,-150487,
    -150172,-149859,-149546,-149235,-148924,-148615,-148307,-148000,
    -147693,-147388,-147084,-146782,-146480,-146179,-145879,-145580,
    -145282,-144986,-144690,-144395,-144101,-143808,-143517,-143226,
    -142936,-142647,-142359,-142072,-141786,-141501,-141217,-140934,
    -140651,-140370,-140090,-139810,-139532,-139254,-138977,-138701,
    -138426,-138152,-137879,-137607,-137335,-137065,-136795,-136526,
    -136258,-135991,-135725,-135459,-135195,-134931,-134668,-134406,
    -134145,-133884,-133625,-133366,-133108,-132851,-132594,-132339,
    -132084,-131830,-131576,-131324,-131072,-130821,-130571,-130322,
    -130073,-129825,-129578,-129332,-129086,-128841,-128597,-128353,
    -128111,-127869,-127627,-127387,-127147,-126908,-126669,-126432,
    -126195,-125959,-125723,-125488,-125254,-125020,-124787,-124555,
    -124324,-124093,-123863,-123633,-123404,-123176,-122949,-122722,
    -122496,-122270,-122045,-121821,-121597,-121374,-121152,-120930,
    -120709,-120489,-120269,-120050,-119831,-119613,-119396,-119179,
    -118963,-118747,-118532,-118318,-118104,-117891,-117678,-117466,
    -117254,-117044,-116833,-116623,-116414,-116206,-115998,-115790,
    -115583,-115377,-115171,-114966,-114761,-114557,-114354,-114151,
    -113948,-113746,-113545,-113344,-113143,-112944,-112744,-112546,
    -112347,-112150,-111952,-111756,-111560,-111364,-111169,-110974,
    -110780,-110586,-110393,-110200,-110008,-109817,-109626,-109435,
    -109245,-109055,-108866,-108677,-108489,-108301,-108114,-107927,
    -107741,-107555,-107369,-107184,-107000,-106816,-106632,-106449,
    -106266,-106084,-105902,-105721,-105540,-105360,-105180,-105000,
    -104821,-104643,-104465,-104287,-104109,-103933,-103756,-103580,
    -103404,-103229,-103054,-102880,-102706,-102533,-102360,-102187,
    -102015,-101843,-101671,-101500,-101330,-101159,-100990,-100820,
    -100651,-100482,-100314,-100146,-99979,-99812,-99645,-99479,
    -99313,-99148,-98982,-98818,-98653,-98489,-98326,-98163,
    -98000,-97837,-97675,-97513,-97352,-97191,-97030,-96870,
    -96710,-96551,-96391,-96233,-96074,-95916,-95758,-95601,
    -95444,-95287,-95131,-94975,-94819,-94664,-94509,-94354,
    -94200,-94046,-93892,-93739,-93586,-93434,-93281,-93129,
    -92978,-92826,-92675,-92525,-92375,-92225,-92075,-91926,
    -91777,-91628,-91480,-91332,-91184,-91036,-90889,-90742,
    -90596,-90450,-90304,-90158,-90013,-89868,-89724,-89579,
    -89435,-89292,-89148,-89005,-88862,-88720,-88577,-88435,
    -88294,-88152,-88011,-87871,-87730,-87590,-87450,-87310,
    -87171,-87032,-86893,-86755,-86616,-86479,-86341,-86204,
    -86066,-85930,-85793,-85657,-85521,-85385,-85250,-85114,
    -84980,-84845,-84710,-84576,-84443,-84309,-84176,-84043,
    -83910,-83777,-83645,-83513,-83381,-83250,-83118,-82987,
    -82857,-82726,-82596,-82466,-82336,-82207,-82078,-81949,
    -81820,-81691,-81563,-81435,-81307,-81180,-81053,-80925,
    -80799,-80672,-80546,-80420,-80294,-80168,-80043,-79918,
    -79793,-79668,-79544,-79420,-79296,-79172,-79048,-78925,
    -78802,-78679,-78557,-78434,-78312,-78190,-78068,-77947,
    -77826,-77705,-77584,-77463,-77343,-77223,-77103,-76983,
    -76864,-76744,-76625,-76506,-76388,-76269,-76151,-76033,
    -75915,-75797,-75680,-75563,-75446,-75329,-75213,-75096,
    -74980,-74864,-74748,-74633,-74517,-74402,-74287,-74172,
    -74058,-73944,-73829,-73715,-73602,-73488,-73375,-73262,
    -73149,-73036,-72923,-72811,-72699,-72587,-72475,-72363,
    -72252,-72140,-72029,-71918,-71808,-71697,-71587,-71477,
    -71367,-71257,-71147,-71038,-70929,-70820,-70711,-70602,
    -70494,-70385,-70277,-70169,-70061,-69954,-69846,-69739,
    -69632,-69525,-69418,-69312,-69205,-69099,-68993,-68887,
    -68781,-68676,-68570,-68465,-68360,-68255,-68151,-68046,
    -67942,-67837,-67733,-67629,-67526,-67422,-67319,-67216,
    -67113,-67010,-66907,-66804,-66702,-66600,-66498,-66396,
    -66294,-66192,-66091,-65989,-65888,-65787,-65686,-65586,
    -65485,-65385,-65285,-65185,-65085,-64985,-64885,-64786,
    -64687,-64587,-64488,-64389,-64291,-64192,-64094,-63996,
    -63897,-63799,-63702,-63604,-63506,-63409,-63312,-63215,
    -63118,-63021,-62924,-62828,-62731,-62635,-62539,-62443,
    -62347,-62251,-62156,-62060,-61965,-61870,-61775,-61680,
    -61585,-61491,-61396,-61302,-61208,-61114,-61020,-60926,
    -60833,-60739,-60646,-60552,-60459,-60366,-60273,-60181,
    -60088,-59996,-59903,-59811,-59719,-59627,-59535,-59444,
    -59352,-59261,-59169,-59078,-58987,-58896,-58805,-58715,
    -58624,-58534,-58443,-58353,-58263,-58173,-58083,-57994,
    -57904,-57815,-57725,-57636,-57547,-57458,-57369,-57281,
    -57192,-57104,-57015,-56927,-56839,-56751,-56663,-56575,
    -56487,-56400,-56312,-56225,-56138,-56051,-55964,-55877,
    -55790,-55704,-55617,-55531,-55444,-55358,-55272,-55186,
    -55100,-55015,-54929,-54843,-54758,-54673,-54587,-54502,
    -54417,-54333,-54248,-54163,-54079,-53994,-53910,-53826,
    -53741,-53657,-53574,-53490,-53406,-53322,-53239,-53156,
    -53072,-52989,-52906,-52823,-52740,-52657,-52575,-52492,
    -52410,-52327,-52245,-52163,-52081,-51999,-51917,-51835,
    -51754,-51672,-51591,-51509,-51428,-51347,-51266,-51185,
    -51104,-51023,-50942,-50862,-50781,-50701,-50621,-50540,
    -50460,-50380,-50300,-50221,-50141,-50061,-49982,-49902,
    -49823,-49744,-49664,-49585,-49506,-49427,-49349,-49270,
    -49191,-49113,-49034,-48956,-48878,-48799,-48721,-48643,
    -48565,-48488,-48410,-48332,-48255,-48177,-48100,-48022,
    -47945,-47868,-47791,-47714,-47637,-47560,-47484,-47407,
    -47331,-47254,-47178,-47102,-47025,-46949,-46873,-46797,
    -46721,-46646,-46570,-46494,-46419,-46343,-46268,-46193,
    -46118,-46042,-45967,-45892,-45818,-45743,-45668,-45593,
    -45519,-45444,-45370,-45296,-45221,-45147,-45073,-44999,
    -44925,-44851,-44778,-44704,-44630,-44557,-44483,-44410,
    -44337,-44263,-44190,-44117,-44044,-43971,-43898,-43826,
    -43753,-43680,-43608,-43535,-43463,-43390,-43318,-43246,
    -43174,-43102,-43030,-42958,-42886,-42814,-42743,-42671,
    -42600,-42528,-42457,-42385,-42314,-42243,-42172,-42101,
    -42030,-41959,-41888,-41817,-41747,-41676,-41605,-41535,
    -41465,-41394,-41324,-41254,-41184,-41113,-41043,-40973,
    -40904,-40834,-40764,-40694,-40625,-40555,-40486,-40416,
    -40347,-40278,-40208,-40139,-40070,-40001,-39932,-39863,
    -39794,-39726,-39657,-39588,-39520,-39451,-39383,-39314,
    -39246,-39178,-39110,-39042,-38973,-38905,-38837,-38770,
    -38702,-38634,-38566,-38499,-38431,-38364,-38296,-38229,
    -38161,-38094,-38027,-37960,-37893,-37826,-37759,-37692,
    -37625,-37558,-37491,-37425,-37358,-37291,-37225,-37158,
    -37092,-37026,-36959,-36893,-36827,-36761,-36695,-36629,
    -36563,-36497,-36431,-36365,-36300,-36234,-36168,-36103,
    -36037,-35972,-35907,-35841,-35776,-35711,-35646,-35580,
    -35515,-35450,-35385,-35321,-35256,-35191,-35126,-35062,
    -34997,-34932,-34868,-34803,-34739,-34675,-34610,-34546,
    -34482,-34418,-34354,-34289,-34225,-34162,-34098,-34034,
    -33970,-33906,-33843,-33779,-33715,-33652,-33588,-33525,
    -33461,-33398,-33335,-33272,-33208,-33145,-33082,-33019,
    -32956,-32893,-32830,-32767,-32705,-32642,-32579,-32516,
    -32454,-32391,-32329,-32266,-32204,-32141,-32079,-32017,
    -31955,-31892,-31830,-31768,-31706,-31644,-31582,-31520,
    -31458,-31396,-31335,-31273,-31211,-31150,-31088,-31026,
    -30965,-30904,-30842,-30781,-30719,-30658,-30597,-30536,
    -30474,-30413,-30352,-30291,-30230,-30169,-30108,-30048,
    -29987,-29926,-29865,-29805,-29744,-29683,-29623,-29562,
    -29502,-29441,-29381,-29321,-29260,-29200,-29140,-29080,
    -29020,-28959,-28899,-28839,-28779,-28719,-28660,-28600,
    -28540,-28480,-28420,-28361,-28301,-28241,-28182,-28122,
    -28063,-28003,-27944,-27884,-27825,-27766,-27707,-27647,
    -27588,-27529,-27470,-27411,-27352,-27293,-27234,-27175,
    -27116,-27057,-26998,-26940,-26881,-26822,-26763,-26705,
    -26646,-26588,-26529,-26471,-26412,-26354,-26295,-26237,
    -26179,-26120,-26062,-26004,-25946,-25888,-25830,-25772,
    -25714,-25656,-25598,-25540,-25482,-25424,-25366,-25308,
    -25251,-25193,-25135,-25078,-25020,-24962,-24905,-24847,
    -24790,-24732,-24675,-24618,-24560,-24503,-24446,-24389,
    -24331,-24274,-24217,-24160,-24103,-24046,-23989,-23932,
    -23875,-23818,-23761,-23704,-23647,-23591,-23534,-23477,
    -23420,-23364,-23307,-23250,-23194,-23137,-23081,-23024,
    -22968,-22911,-22855,-22799,-22742,-22686,-22630,-22573,
    -22517,-22461,-22405,-22349,-22293,-22237,-22181,-22125,
    -22069,-22013,-21957,-21901,-21845,-21789,-21733,-21678,
    -21622,-21566,-21510,-21455,-21399,-21343,-21288,-21232,
    -21177,-21121,-21066,-21010,-20955,-20900,-20844,-20789,
    -20734,-20678,-20623,-20568,-20513,-20457,-20402,-20347,
    -20292,-20237,-20182,-20127,-20072,-20017,-19962,-19907,
    -19852,-19797,-19742,-19688,-19633,-19578,-19523,-19469,
    -19414,-19359,-19305,-19250,-19195,-19141,-19086,-19032,
    -18977,-18923,-18868,-18814,-18760,-18705,-18651,-18597,
    -18542,-18488,-18434,-18380,-18325,-18271,-18217,-18163,
    -18109,-18055,-18001,-17946,-17892,-17838,-17784,-17731,
    -17677,-17623,-17569,-17515,-17461,-17407,-17353,-17300,
    -17246,-17192,-17138,-17085,-17031,-16977,-16924,-16870,
    -16817,-16763,-16710,-16656,-16603,-16549,-16496,-16442,
    -16389,-16335,-16282,-16229,-16175,-16122,-16069,-16015,
    -15962,-15909,-15856,-15802,-15749,-15696,-15643,-15590,
    -15537,-15484,-15431,-15378,-15325,-15272,-15219,-15166,
    -15113,-15060,-15007,-14954,-14901,-14848,-14795,-14743,
    -14690,-14637,-14584,-14531,-14479,-14426,-14373,-14321,
    -14268,-14215,-14163,-14110,-14057,-14005,-13952,-13900,
    -13847,-13795,-13742,-13690,-13637,-13585,-13533,-13480,
    -13428,-13375,-13323,-13271,-13218,-13166,-13114,-13062,
    -13009,-12957,-12905,-12853,-12800,-12748,-12696,-12644,
    -12592,-12540,-12488,-12436,-12383,-12331,-12279,-12227,
    -12175,-12123,-12071,-12019,-11967,-11916,-11864,-11812,
    -11760,-11708,-11656,-11604,-11552,-11501,-11449,-11397,
    -11345,-11293,-11242,-11190,-11138,-11086,-11035,-10983,
    -10931,-10880,-10828,-10777,-10725,-10673,-10622,-10570,
    -10519,-10467,-10415,-10364,-10312,-10261,-10209,-10158,
    -10106,-10055,-10004,-9952,-9901,-9849,-9798,-9747,
    -9695,-9644,-9592,-9541,-9490,-9438,-9387,-9336,
    -9285,-9233,-9182,-9131,-9080,-9028,-8977,-8926,
    -8875,-8824,-8772,-8721,-8670,-8619,-8568,-8517,
    -8466,-8414,-8363,-8312,-8261,-8210,-8159,-8108,
    -8057,-8006,-7955,-7904,-7853,-7802,-7751,-7700,
    -7649,-7598,-7547,-7496,-7445,-7395,-7344,-7293,
    -7242,-7191,-7140,-7089,-7038,-6988,-6937,-6886,
    -6835,-6784,-6733,-6683,-6632,-6581,-6530,-6480,
    -6429,-6378,-6327,-6277,-6226,-6175,-6124,-6074,
    -6023,-5972,-5922,-5871,-5820,-5770,-5719,-5668,
    -5618,-5567,-5517,-5466,-5415,-5365,-5314,-5264,
    -5213,-5162,-5112,-5061,-5011,-4960,-4910,-4859,
    -4808,-4758,-4707,-4657,-4606,-4556,-4505,-4455,
    -4404,-4354,-4303,-4253,-4202,-4152,-4101,-4051,
    -4001,-3950,-3900,-3849,-3799,-3748,-3698,-3648,
    -3597,-3547,-3496,-3446,-3395,-3345,-3295,-3244,
    -3194,-3144,-3093,-3043,-2992,-2942,-2892,-2841,
    -2791,-2741,-2690,-2640,-2590,-2539,-2489,-2439,
    -2388,-2338,-2288,-2237,-2187,-2137,-2086,-2036,
    -1986,-1935,-1885,-1835,-1784,-1734,-1684,-1633,
    -1583,-1533,-1483,-1432,-1382,-1332,-1281,-1231,
    -1181,-1131,-1080,-1030,-980,-929,-879,-829,
    -779,-728,-678,-628,-578,-527,-477,-427,
    -376,-326,-276,-226,-175,-125,-75,-25,
    25,75,125,175,226,276,326,376,
    427,477,527,578,628,678,728,779,
    829,879,929,980,1030,1080,1131,1181,
    1231,1281,1332,1382,1432,1483,1533,1583,
    1633,1684,1734,1784,1835,1885,1935,1986,
    2036,2086,2137,2187,2237,2288,2338,2388,
    2439,2489,2539,2590,2640,2690,2741,2791,
    2841,2892,2942,2992,3043,3093,3144,3194,
    3244,3295,3345,3395,3446,3496,3547,3597,
    3648,3698,3748,3799,3849,3900,3950,4001,
    4051,4101,4152,4202,4253,4303,4354,4404,
    4455,4505,4556,4606,4657,4707,4758,4808,
    4859,4910,4960,5011,5061,5112,5162,5213,
    5264,5314,5365,5415,5466,5517,5567,5618,
    5668,5719,5770,5820,5871,5922,5972,6023,
    6074,6124,6175,6226,6277,6327,6378,6429,
    6480,6530,6581,6632,6683,6733,6784,6835,
    6886,6937,6988,7038,7089,7140,7191,7242,
    7293,7344,7395,7445,7496,7547,7598,7649,
    7700,7751,7802,7853,7904,7955,8006,8057,
    8108,8159,8210,8261,8312,8363,8414,8466,
    8517,8568,8619,8670,8721,8772,8824,8875,
    8926,8977,9028,9080,9131,9182,9233,9285,
    9336,9387,9438,9490,9541,9592,9644,9695,
    9747,9798,9849,9901,9952,10004,10055,10106,
    10158,10209,10261,10312,10364,10415,10467,10519,
    10570,10622,10673,10725,10777,10828,10880,10931,
    10983,11035,11086,11138,11190,11242,11293,11345,
    11397,11449,11501,11552,11604,11656,11708,11760,
    11812,11864,11916,11967,12019,12071,12123,12175,
    12227,12279,12331,12383,12436,12488,12540,12592,
    12644,12696,12748,12800,12853,12905,12957,13009,
    13062,13114,13166,13218,13271,13323,13375,13428,
    13480,13533,13585,13637,13690,13742,13795,13847,
    13900,13952,14005,14057,14110,14163,14215,14268,
    14321,14373,14426,14479,14531,14584,14637,14690,
    14743,14795,14848,14901,14954,15007,15060,15113,
    15166,15219,15272,15325,15378,15431,15484,15537,
    15590,15643,15696,15749,15802,15856,15909,15962,
    16015,16069,16122,16175,16229,16282,16335,16389,
    16442,16496,16549,16603,16656,16710,16763,16817,
    16870,16924,16977,17031,17085,17138,17192,17246,
    17300,17353,17407,17461,17515,17569,17623,17677,
    17731,17784,17838,17892,17946,18001,18055,18109,
    18163,18217,18271,18325,18380,18434,18488,18542,
    18597,18651,18705,18760,18814,18868,18923,18977,
    19032,19086,19141,19195,19250,19305,19359,19414,
    19469,19523,19578,19633,19688,19742,19797,19852,
    19907,19962,20017,20072,20127,20182,20237,20292,
    20347,20402,20457,20513,20568,20623,20678,20734,
    20789,20844,20900,20955,21010,21066,21121,21177,
    21232,21288,21343,21399,21455,21510,21566,21622,
    21678,21733,21789,21845,21901,21957,22013,22069,
    22125,22181,22237,22293,22349,22405,22461,22517,
    22573,22630,22686,22742,22799,22855,22911,22968,
    23024,23081,23137,23194,23250,23307,23364,23420,
    23477,23534,23591,23647,23704,23761,23818,23875,
    23932,23989,24046,24103,24160,24217,24274,24331,
    24389,24446,24503,24560,24618,24675,24732,24790,
    24847,24905,24962,25020,25078,25135,25193,25251,
    25308,25366,25424,25482,25540,25598,25656,25714,
    25772,25830,25888,25946,26004,26062,26120,26179,
    26237,26295,26354,26412,26471,26529,26588,26646,
    26705,26763,26822,26881,26940,26998,27057,27116,
    27175,27234,27293,27352,27411,27470,27529,27588,
    27647,27707,27766,27825,27884,27944,28003,28063,
    28122,28182,28241,28301,28361,28420,28480,28540,
    28600,28660,28719,28779,28839,28899,28959,29020,
    29080,29140,29200,29260,29321,29381,29441,29502,
    29562,29623,29683,29744,29805,29865,29926,29987,
    30048,30108,30169,30230,30291,30352,30413,30474,
    30536,30597,30658,30719,30781,30842,30904,30965,
    31026,31088,31150,31211,31273,31335,31396,31458,
    31520,31582,31644,31706,31768,31830,31892,31955,
    32017,32079,32141,32204,32266,32329,32391,32454,
    32516,32579,32642,32705,32767,32830,32893,32956,
    33019,33082,33145,33208,33272,33335,33398,33461,
    33525,33588,33652,33715,33779,33843,33906,33970,
    34034,34098,34162,34225,34289,34354,34418,34482,
    34546,34610,34675,34739,34803,34868,34932,34997,
    35062,35126,35191,35256,35321,35385,35450,35515,
    35580,35646,35711,35776,35841,35907,35972,36037,
    36103,36168,36234,36300,36365,36431,36497,36563,
    36629,36695,36761,36827,36893,36959,37026,37092,
    37158,37225,37291,37358,37425,37491,37558,37625,
    37692,37759,37826,37893,37960,38027,38094,38161,
    38229,38296,38364,38431,38499,38566,38634,38702,
    38770,38837,38905,38973,39042,39110,39178,39246,
    39314,39383,39451,39520,39588,39657,39726,39794,
    39863,39932,40001,40070,40139,40208,40278,40347,
    40416,40486,40555,40625,40694,40764,40834,40904,
    40973,41043,41113,41184,41254,41324,41394,41465,
    41535,41605,41676,41747,41817,41888,41959,42030,
    42101,42172,42243,42314,42385,42457,42528,42600,
    42671,42743,42814,42886,42958,43030,43102,43174,
    43246,43318,43390,43463,43535,43608,43680,43753,
    43826,43898,43971,44044,44117,44190,44263,44337,
    44410,44483,44557,44630,44704,44778,44851,44925,
    44999,45073,45147,45221,45296,45370,45444,45519,
    45593,45668,45743,45818,45892,45967,46042,46118,
    46193,46268,46343,46419,46494,46570,46646,46721,
    46797,46873,46949,47025,47102,47178,47254,47331,
    47407,47484,47560,47637,47714,47791,47868,47945,
    48022,48100,48177,48255,48332,48410,48488,48565,
    48643,48721,48799,48878,48956,49034,49113,49191,
    49270,49349,49427,49506,49585,49664,49744,49823,
    49902,49982,50061,50141,50221,50300,50380,50460,
    50540,50621,50701,50781,50862,50942,51023,51104,
    51185,51266,51347,51428,51509,51591,51672,51754,
    51835,51917,51999,52081,52163,52245,52327,52410,
    52492,52575,52657,52740,52823,52906,52989,53072,
    53156,53239,53322,53406,53490,53574,53657,53741,
    53826,53910,53994,54079,54163,54248,54333,54417,
    54502,54587,54673,54758,54843,54929,55015,55100,
    55186,55272,55358,55444,55531,55617,55704,55790,
    55877,55964,56051,56138,56225,56312,56400,56487,
    56575,56663,56751,56839,56927,57015,57104,57192,
    57281,57369,57458,57547,57636,57725,57815,57904,
    57994,58083,58173,58263,58353,58443,58534,58624,
    58715,58805,58896,58987,59078,59169,59261,59352,
    59444,59535,59627,59719,59811,59903,59996,60088,
    60181,60273,60366,60459,60552,60646,60739,60833,
    60926,61020,61114,61208,61302,61396,61491,61585,
    61680,61775,61870,61965,62060,62156,62251,62347,
    62443,62539,62635,62731,62828,62924,63021,63118,
    63215,63312,63409,63506,63604,63702,63799,63897,
    63996,64094,64192,64291,64389,64488,64587,64687,
    64786,64885,64985,65085,65185,65285,65385,65485,
    65586,65686,65787,65888,65989,66091,66192,66294,
    66396,66498,66600,66702,66804,66907,67010,67113,
    67216,67319,67422,67526,67629,67733,67837,67942,
    68046,68151,68255,68360,68465,68570,68676,68781,
    68887,68993,69099,69205,69312,69418,69525,69632,
    69739,69846,69954,70061,70169,70277,70385,70494,
    70602,70711,70820,70929,71038,71147,71257,71367,
    71477,71587,71697,71808,71918,72029,72140,72252,
    72363,72475,72587,72699,72811,72923,73036,73149,
    73262,73375,73488,73602,73715,73829,73944,74058,
    74172,74287,74402,74517,74633,74748,74864,74980,
    75096,75213,75329,75446,75563,75680,75797,75915,
    76033,76151,76269,76388,76506,76625,76744,76864,
    76983,77103,77223,77343,77463,77584,77705,77826,
    77947,78068,78190,78312,78434,78557,78679,78802,
    78925,79048,79172,79296,79420,79544,79668,79793,
    79918,80043,80168,80294,80420,80546,80672,80799,
    80925,81053,81180,81307,81435,81563,81691,81820,
    81949,82078,82207,82336,82466,82596,82726,82857,
    82987,83118,83250,83381,83513,83645,83777,83910,
    84043,84176,84309,84443,84576,84710,84845,84980,
    85114,85250,85385,85521,85657,85793,85930,86066,
    86204,86341,86479,86616,86755,86893,87032,87171,
    87310,87450,87590,87730,87871,88011,88152,88294,
    88435,88577,88720,88862,89005,89148,89292,89435,
    89579,89724,89868,90013,90158,90304,90450,90596,
    90742,90889,91036,91184,91332,91480,91628,91777,
    91926,92075,92225,92375,92525,92675,92826,92978,
    93129,93281,93434,93586,93739,93892,94046,94200,
    94354,94509,94664,94819,94975,95131,95287,95444,
    95601,95758,95916,96074,96233,96391,96551,96710,
    96870,97030,97191,97352,97513,97675,97837,98000,
    98163,98326,98489,98653,98818,98982,99148,99313,
    99479,99645,99812,99979,100146,100314,100482,100651,
    100820,100990,101159,101330,101500,101671,101843,102015,
    102187,102360,102533,102706,102880,103054,103229,103404,
    103580,103756,103933,104109,104287,104465,104643,104821,
    105000,105180,105360,105540,105721,105902,106084,106266,
    106449,106632,106816,107000,107184,107369,107555,107741,
    107927,108114,108301,108489,108677,108866,109055,109245,
    109435,109626,109817,110008,110200,110393,110586,110780,
    110974,111169,111364,111560,111756,111952,112150,112347,
    112546,112744,112944,113143,113344,113545,113746,113948,
    114151,114354,114557,114761,114966,115171,115377,115583,
    115790,115998,116206,116414,116623,116833,117044,117254,
    117466,117678,117891,118104,118318,118532,118747,118963,
    119179,119396,119613,119831,120050,120269,120489,120709,
    120930,121152,121374,121597,121821,122045,122270,122496,
    122722,122949,123176,123404,123633,123863,124093,124324,
    124555,124787,125020,125254,125488,125723,125959,126195,
    126432,126669,126908,127147,127387,127627,127869,128111,
    128353,128597,128841,129086,129332,129578,129825,130073,
    130322,130571,130821,131072,131324,131576,131830,132084,
    132339,132594,132851,133108,133366,133625,133884,134145,
    134406,134668,134931,135195,135459,135725,135991,136258,
    136526,136795,137065,137335,137607,137879,138152,138426,
    138701,138977,139254,139532,139810,140090,140370,140651,
    140934,141217,141501,141786,142072,142359,142647,142936,
    143226,143517,143808,144101,144395,144690,144986,145282,
    145580,145879,146179,146480,146782,147084,147388,147693,
    148000,148307,148615,148924,149235,149546,149859,150172,
    150487,150803,151120,151438,151757,152077,152399,152722,
    153045,153370,153697,154024,154352,154682,155013,155345,
    155678,156013,156349,156686,157024,157363,157704,158046,
    158389,158734,159079,159427,159775,160125,160476,160828,
    161182,161537,161893,162251,162610,162970,163332,163695,
    164060,164426,164793,165162,165532,165904,166277,166651,
    167027,167405,167784,168164,168546,168930,169315,169701,
    170089,170479,170870,171263,171657,172053,172451,172850,
    173251,173653,174057,174463,174870,175279,175690,176102,
    176516,176932,177349,177769,178190,178612,179037,179463,
    179891,180321,180753,181186,181622,182059,182498,182939,
    183382,183827,184274,184722,185173,185625,186080,186536,
    186995,187455,187918,188382,188849,189318,189789,190261,
    190736,191213,191693,192174,192658,193143,193631,194122,
    194614,195109,195606,196105,196606,197110,197616,198125,
    198636,199149,199664,200182,200703,201226,201751,202279,
    202809,203342,203878,204416,204956,205500,206045,206594,
    207145,207699,208255,208815,209376,209941,210509,211079,
    211652,212228,212807,213389,213973,214561,215151,215745,
    216341,216941,217544,218149,218758,219370,219985,220603,
    221225,221849,222477,223108,223743,224381,225022,225666,
    226314,226966,227621,228279,228941,229606,230275,230948,
    231624,232304,232988,233676,234367,235062,235761,236463,
    237170,237881,238595,239314,240036,240763,241493,242228,
    242967,243711,244458,245210,245966,246727,247492,248261,
    249035,249813,250596,251384,252176,252973,253774,254581,
    255392,256208,257029,257855,258686,259522,260363,261209,
    262060,262917,263779,264646,265519,266397,267280,268169,
    269064,269965,270871,271782,272700,273624,274553,275489,
    276430,277378,278332,279292,280258,281231,282210,283195,
    284188,285186,286192,287204,288223,289249,290282,291322,
    292369,293423,294485,295554,296630,297714,298805,299904,
    301011,302126,303248,304379,305517,306664,307819,308983,
    310154,311335,312524,313721,314928,316143,317368,318601,
    319844,321097,322358,323629,324910,326201,327502,328812,
    330133,331464,332805,334157,335519,336892,338276,339671,
    341078,342495,343924,345364,346816,348280,349756,351244,
    352744,354257,355783,357321,358872,360436,362013,363604,
    365208,366826,368459,370105,371765,373440,375130,376835,
    378555,380290,382040,383807,385589,387387,389202,391034,
    392882,394747,396630,398530,400448,402384,404338,406311,
    408303,410314,412344,414395,416465,418555,420666,422798,
    424951,427125,429321,431540,433781,436045,438332,440643,
    442978,445337,447720,450129,452564,455024,457511,460024,
    462565,465133,467730,470355,473009,475692,478406,481150,
    483925,486732,489571,492443,495348,498287,501261,504269,
    507313,510394,513512,516667,519861,523094,526366,529680,
    533034,536431,539870,543354,546881,550455,554074,557741,
    561456,565221,569035,572901,576818,580789,584815,588896,
    593033,597229,601483,605798,610174,614613,619117,623686,
    628323,633028,637803,642651,647572,652568,657640,662792,
    668024,673338,678737,684223,689797,695462,701219,707072,
    713023,719074,725227,731486,737853,744331,750922,757631,
    764460,771411,778490,785699,793041,800521,808143,815910,
    823827,831898,840127,848520,857081,865817,874730,883829,
    893117,902602,912289,922186,932298,942633,953199,964003,
    975054,986361,997931,1009774,1021901,1034322,1047046,1060087,
    1073455,1087164,1101225,1115654,1130465,1145673,1161294,1177345,
    1193846,1210813,1228269,1246234,1264730,1283783,1303416,1323658,
    1344537,1366084,1388330,1411312,1435065,1459630,1485049,1511367,
    1538632,1566898,1596220,1626658,1658278,1691149,1725348,1760956,
    1798063,1836758,1877161,1919378,1963536,2009771,2058233,2109087,
    2162516,2218719,2277919,2340362,2406322,2476104,2550052,2628549,
    2712030,2800983,2895966,2997613,3106651,3223918,3350381,3487165,
    3635590,3797206,3973855,4167737,4381502,4618375,4882318,5178251,
    5512368,5892567,6329090,6835455,7429880,8137527,8994149,10052327,
    11392683,13145455,15535599,18988036,24413316,34178904,56965752,170910304
)]!

const finesine = [i32(
25,75,125,175,226,276,326,376,
    427,477,527,578,628,678,728,779,
    829,879,929,980,1030,1080,1130,1181,
    1231,1281,1331,1382,1432,1482,1532,1583,
    1633,1683,1733,1784,1834,1884,1934,1985,
    2035,2085,2135,2186,2236,2286,2336,2387,
    2437,2487,2537,2587,2638,2688,2738,2788,
    2839,2889,2939,2989,3039,3090,3140,3190,
    3240,3291,3341,3391,3441,3491,3541,3592,
    3642,3692,3742,3792,3843,3893,3943,3993,
    4043,4093,4144,4194,4244,4294,4344,4394,
    4445,4495,4545,4595,4645,4695,4745,4796,
    4846,4896,4946,4996,5046,5096,5146,5197,
    5247,5297,5347,5397,5447,5497,5547,5597,
    5647,5697,5748,5798,5848,5898,5948,5998,
    6048,6098,6148,6198,6248,6298,6348,6398,
    6448,6498,6548,6598,6648,6698,6748,6798,
    6848,6898,6948,6998,7048,7098,7148,7198,
    7248,7298,7348,7398,7448,7498,7548,7598,
    7648,7697,7747,7797,7847,7897,7947,7997,
    8047,8097,8147,8196,8246,8296,8346,8396,
    8446,8496,8545,8595,8645,8695,8745,8794,
    8844,8894,8944,8994,9043,9093,9143,9193,
    9243,9292,9342,9392,9442,9491,9541,9591,
    9640,9690,9740,9790,9839,9889,9939,9988,
    10038,10088,10137,10187,10237,10286,10336,10386,
    10435,10485,10534,10584,10634,10683,10733,10782,
    10832,10882,10931,10981,11030,11080,11129,11179,
    11228,11278,11327,11377,11426,11476,11525,11575,
    11624,11674,11723,11773,11822,11872,11921,11970,
    12020,12069,12119,12168,12218,12267,12316,12366,
    12415,12464,12514,12563,12612,12662,12711,12760,
    12810,12859,12908,12957,13007,13056,13105,13154,
    13204,13253,13302,13351,13401,13450,13499,13548,
    13597,13647,13696,13745,13794,13843,13892,13941,
    13990,14040,14089,14138,14187,14236,14285,14334,
    14383,14432,14481,14530,14579,14628,14677,14726,
    14775,14824,14873,14922,14971,15020,15069,15118,
    15167,15215,15264,15313,15362,15411,15460,15509,
    15557,15606,15655,15704,15753,15802,15850,15899,
    15948,15997,16045,16094,16143,16191,16240,16289,
    16338,16386,16435,16484,16532,16581,16629,16678,
    16727,16775,16824,16872,16921,16970,17018,17067,
    17115,17164,17212,17261,17309,17358,17406,17455,
    17503,17551,17600,17648,17697,17745,17793,17842,
    17890,17939,17987,18035,18084,18132,18180,18228,
    18277,18325,18373,18421,18470,18518,18566,18614,
    18663,18711,18759,18807,18855,18903,18951,19000,
    19048,19096,19144,19192,19240,19288,19336,19384,
    19432,19480,19528,19576,19624,19672,19720,19768,
    19816,19864,19912,19959,20007,20055,20103,20151,
    20199,20246,20294,20342,20390,20438,20485,20533,
    20581,20629,20676,20724,20772,20819,20867,20915,
    20962,21010,21057,21105,21153,21200,21248,21295,
    21343,21390,21438,21485,21533,21580,21628,21675,
    21723,21770,21817,21865,21912,21960,22007,22054,
    22102,22149,22196,22243,22291,22338,22385,22433,
    22480,22527,22574,22621,22668,22716,22763,22810,
    22857,22904,22951,22998,23045,23092,23139,23186,
    23233,23280,23327,23374,23421,23468,23515,23562,
    23609,23656,23703,23750,23796,23843,23890,23937,
    23984,24030,24077,24124,24171,24217,24264,24311,
    24357,24404,24451,24497,24544,24591,24637,24684,
    24730,24777,24823,24870,24916,24963,25009,25056,
    25102,25149,25195,25241,25288,25334,25381,25427,
    25473,25520,25566,25612,25658,25705,25751,25797,
    25843,25889,25936,25982,26028,26074,26120,26166,
    26212,26258,26304,26350,26396,26442,26488,26534,
    26580,26626,26672,26718,26764,26810,26856,26902,
    26947,26993,27039,27085,27131,27176,27222,27268,
    27313,27359,27405,27450,27496,27542,27587,27633,
    27678,27724,27770,27815,27861,27906,27952,27997,
    28042,28088,28133,28179,28224,28269,28315,28360,
    28405,28451,28496,28541,28586,28632,28677,28722,
    28767,28812,28858,28903,28948,28993,29038,29083,
    29128,29173,29218,29263,29308,29353,29398,29443,
    29488,29533,29577,29622,29667,29712,29757,29801,
    29846,29891,29936,29980,30025,30070,30114,30159,
    30204,30248,30293,30337,30382,30426,30471,30515,
    30560,30604,30649,30693,30738,30782,30826,30871,
    30915,30959,31004,31048,31092,31136,31181,31225,
    31269,31313,31357,31402,31446,31490,31534,31578,
    31622,31666,31710,31754,31798,31842,31886,31930,
    31974,32017,32061,32105,32149,32193,32236,32280,
    32324,32368,32411,32455,32499,32542,32586,32630,
    32673,32717,32760,32804,32847,32891,32934,32978,
    33021,33065,33108,33151,33195,33238,33281,33325,
    33368,33411,33454,33498,33541,33584,33627,33670,
    33713,33756,33799,33843,33886,33929,33972,34015,
    34057,34100,34143,34186,34229,34272,34315,34358,
    34400,34443,34486,34529,34571,34614,34657,34699,
    34742,34785,34827,34870,34912,34955,34997,35040,
    35082,35125,35167,35210,35252,35294,35337,35379,
    35421,35464,35506,35548,35590,35633,35675,35717,
    35759,35801,35843,35885,35927,35969,36011,36053,
    36095,36137,36179,36221,36263,36305,36347,36388,
    36430,36472,36514,36555,36597,36639,36681,36722,
    36764,36805,36847,36889,36930,36972,37013,37055,
    37096,37137,37179,37220,37262,37303,37344,37386,
    37427,37468,37509,37551,37592,37633,37674,37715,
    37756,37797,37838,37879,37920,37961,38002,38043,
    38084,38125,38166,38207,38248,38288,38329,38370,
    38411,38451,38492,38533,38573,38614,38655,38695,
    38736,38776,38817,38857,38898,38938,38979,39019,
    39059,39100,39140,39180,39221,39261,39301,39341,
    39382,39422,39462,39502,39542,39582,39622,39662,
    39702,39742,39782,39822,39862,39902,39942,39982,
    40021,40061,40101,40141,40180,40220,40260,40300,
    40339,40379,40418,40458,40497,40537,40576,40616,
    40655,40695,40734,40773,40813,40852,40891,40931,
    40970,41009,41048,41087,41127,41166,41205,41244,
    41283,41322,41361,41400,41439,41478,41517,41556,
    41595,41633,41672,41711,41750,41788,41827,41866,
    41904,41943,41982,42020,42059,42097,42136,42174,
    42213,42251,42290,42328,42366,42405,42443,42481,
    42520,42558,42596,42634,42672,42711,42749,42787,
    42825,42863,42901,42939,42977,43015,43053,43091,
    43128,43166,43204,43242,43280,43317,43355,43393,
    43430,43468,43506,43543,43581,43618,43656,43693,
    43731,43768,43806,43843,43880,43918,43955,43992,
    44029,44067,44104,44141,44178,44215,44252,44289,
    44326,44363,44400,44437,44474,44511,44548,44585,
    44622,44659,44695,44732,44769,44806,44842,44879,
    44915,44952,44989,45025,45062,45098,45135,45171,
    45207,45244,45280,45316,45353,45389,45425,45462,
    45498,45534,45570,45606,45642,45678,45714,45750,
    45786,45822,45858,45894,45930,45966,46002,46037,
    46073,46109,46145,46180,46216,46252,46287,46323,
    46358,46394,46429,46465,46500,46536,46571,46606,
    46642,46677,46712,46747,46783,46818,46853,46888,
    46923,46958,46993,47028,47063,47098,47133,47168,
    47203,47238,47273,47308,47342,47377,47412,47446,
    47481,47516,47550,47585,47619,47654,47688,47723,
    47757,47792,47826,47860,47895,47929,47963,47998,
    48032,48066,48100,48134,48168,48202,48237,48271,
    48305,48338,48372,48406,48440,48474,48508,48542,
    48575,48609,48643,48676,48710,48744,48777,48811,
    48844,48878,48911,48945,48978,49012,49045,49078,
    49112,49145,49178,49211,49244,49278,49311,49344,
    49377,49410,49443,49476,49509,49542,49575,49608,
    49640,49673,49706,49739,49771,49804,49837,49869,
    49902,49935,49967,50000,50032,50065,50097,50129,
    50162,50194,50226,50259,50291,50323,50355,50387,
    50420,50452,50484,50516,50548,50580,50612,50644,
    50675,50707,50739,50771,50803,50834,50866,50898,
    50929,50961,50993,51024,51056,51087,51119,51150,
    51182,51213,51244,51276,51307,51338,51369,51401,
    51432,51463,51494,51525,51556,51587,51618,51649,
    51680,51711,51742,51773,51803,51834,51865,51896,
    51926,51957,51988,52018,52049,52079,52110,52140,
    52171,52201,52231,52262,52292,52322,52353,52383,
    52413,52443,52473,52503,52534,52564,52594,52624,
    52653,52683,52713,52743,52773,52803,52832,52862,
    52892,52922,52951,52981,53010,53040,53069,53099,
    53128,53158,53187,53216,53246,53275,53304,53334,
    53363,53392,53421,53450,53479,53508,53537,53566,
    53595,53624,53653,53682,53711,53739,53768,53797,
    53826,53854,53883,53911,53940,53969,53997,54026,
    54054,54082,54111,54139,54167,54196,54224,54252,
    54280,54308,54337,54365,54393,54421,54449,54477,
    54505,54533,54560,54588,54616,54644,54672,54699,
    54727,54755,54782,54810,54837,54865,54892,54920,
    54947,54974,55002,55029,55056,55084,55111,55138,
    55165,55192,55219,55246,55274,55300,55327,55354,
    55381,55408,55435,55462,55489,55515,55542,55569,
    55595,55622,55648,55675,55701,55728,55754,55781,
    55807,55833,55860,55886,55912,55938,55965,55991,
    56017,56043,56069,56095,56121,56147,56173,56199,
    56225,56250,56276,56302,56328,56353,56379,56404,
    56430,56456,56481,56507,56532,56557,56583,56608,
    56633,56659,56684,56709,56734,56760,56785,56810,
    56835,56860,56885,56910,56935,56959,56984,57009,
    57034,57059,57083,57108,57133,57157,57182,57206,
    57231,57255,57280,57304,57329,57353,57377,57402,
    57426,57450,57474,57498,57522,57546,57570,57594,
    57618,57642,57666,57690,57714,57738,57762,57785,
    57809,57833,57856,57880,57903,57927,57950,57974,
    57997,58021,58044,58067,58091,58114,58137,58160,
    58183,58207,58230,58253,58276,58299,58322,58345,
    58367,58390,58413,58436,58459,58481,58504,58527,
    58549,58572,58594,58617,58639,58662,58684,58706,
    58729,58751,58773,58795,58818,58840,58862,58884,
    58906,58928,58950,58972,58994,59016,59038,59059,
    59081,59103,59125,59146,59168,59190,59211,59233,
    59254,59276,59297,59318,59340,59361,59382,59404,
    59425,59446,59467,59488,59509,59530,59551,59572,
    59593,59614,59635,59656,59677,59697,59718,59739,
    59759,59780,59801,59821,59842,59862,59883,59903,
    59923,59944,59964,59984,60004,60025,60045,60065,
    60085,60105,60125,60145,60165,60185,60205,60225,
    60244,60264,60284,60304,60323,60343,60363,60382,
    60402,60421,60441,60460,60479,60499,60518,60537,
    60556,60576,60595,60614,60633,60652,60671,60690,
    60709,60728,60747,60766,60785,60803,60822,60841,
    60859,60878,60897,60915,60934,60952,60971,60989,
    61007,61026,61044,61062,61081,61099,61117,61135,
    61153,61171,61189,61207,61225,61243,61261,61279,
    61297,61314,61332,61350,61367,61385,61403,61420,
    61438,61455,61473,61490,61507,61525,61542,61559,
    61577,61594,61611,61628,61645,61662,61679,61696,
    61713,61730,61747,61764,61780,61797,61814,61831,
    61847,61864,61880,61897,61913,61930,61946,61963,
    61979,61995,62012,62028,62044,62060,62076,62092,
    62108,62125,62141,62156,62172,62188,62204,62220,
    62236,62251,62267,62283,62298,62314,62329,62345,
    62360,62376,62391,62407,62422,62437,62453,62468,
    62483,62498,62513,62528,62543,62558,62573,62588,
    62603,62618,62633,62648,62662,62677,62692,62706,
    62721,62735,62750,62764,62779,62793,62808,62822,
    62836,62850,62865,62879,62893,62907,62921,62935,
    62949,62963,62977,62991,63005,63019,63032,63046,
    63060,63074,63087,63101,63114,63128,63141,63155,
    63168,63182,63195,63208,63221,63235,63248,63261,
    63274,63287,63300,63313,63326,63339,63352,63365,
    63378,63390,63403,63416,63429,63441,63454,63466,
    63479,63491,63504,63516,63528,63541,63553,63565,
    63578,63590,63602,63614,63626,63638,63650,63662,
    63674,63686,63698,63709,63721,63733,63745,63756,
    63768,63779,63791,63803,63814,63825,63837,63848,
    63859,63871,63882,63893,63904,63915,63927,63938,
    63949,63960,63971,63981,63992,64003,64014,64025,
    64035,64046,64057,64067,64078,64088,64099,64109,
    64120,64130,64140,64151,64161,64171,64181,64192,
    64202,64212,64222,64232,64242,64252,64261,64271,
    64281,64291,64301,64310,64320,64330,64339,64349,
    64358,64368,64377,64387,64396,64405,64414,64424,
    64433,64442,64451,64460,64469,64478,64487,64496,
    64505,64514,64523,64532,64540,64549,64558,64566,
    64575,64584,64592,64601,64609,64617,64626,64634,
    64642,64651,64659,64667,64675,64683,64691,64699,
    64707,64715,64723,64731,64739,64747,64754,64762,
    64770,64777,64785,64793,64800,64808,64815,64822,
    64830,64837,64844,64852,64859,64866,64873,64880,
    64887,64895,64902,64908,64915,64922,64929,64936,
    64943,64949,64956,64963,64969,64976,64982,64989,
    64995,65002,65008,65015,65021,65027,65033,65040,
    65046,65052,65058,65064,65070,65076,65082,65088,
    65094,65099,65105,65111,65117,65122,65128,65133,
    65139,65144,65150,65155,65161,65166,65171,65177,
    65182,65187,65192,65197,65202,65207,65212,65217,
    65222,65227,65232,65237,65242,65246,65251,65256,
    65260,65265,65270,65274,65279,65283,65287,65292,
    65296,65300,65305,65309,65313,65317,65321,65325,
    65329,65333,65337,65341,65345,65349,65352,65356,
    65360,65363,65367,65371,65374,65378,65381,65385,
    65388,65391,65395,65398,65401,65404,65408,65411,
    65414,65417,65420,65423,65426,65429,65431,65434,
    65437,65440,65442,65445,65448,65450,65453,65455,
    65458,65460,65463,65465,65467,65470,65472,65474,
    65476,65478,65480,65482,65484,65486,65488,65490,
    65492,65494,65496,65497,65499,65501,65502,65504,
    65505,65507,65508,65510,65511,65513,65514,65515,
    65516,65518,65519,65520,65521,65522,65523,65524,
    65525,65526,65527,65527,65528,65529,65530,65530,
    65531,65531,65532,65532,65533,65533,65534,65534,
    65534,65535,65535,65535,65535,65535,65535,65535,
    65535,65535,65535,65535,65535,65535,65535,65534,
    65534,65534,65533,65533,65532,65532,65531,65531,
    65530,65530,65529,65528,65527,65527,65526,65525,
    65524,65523,65522,65521,65520,65519,65518,65516,
    65515,65514,65513,65511,65510,65508,65507,65505,
    65504,65502,65501,65499,65497,65496,65494,65492,
    65490,65488,65486,65484,65482,65480,65478,65476,
    65474,65472,65470,65467,65465,65463,65460,65458,
    65455,65453,65450,65448,65445,65442,65440,65437,
    65434,65431,65429,65426,65423,65420,65417,65414,
    65411,65408,65404,65401,65398,65395,65391,65388,
    65385,65381,65378,65374,65371,65367,65363,65360,
    65356,65352,65349,65345,65341,65337,65333,65329,
    65325,65321,65317,65313,65309,65305,65300,65296,
    65292,65287,65283,65279,65274,65270,65265,65260,
    65256,65251,65246,65242,65237,65232,65227,65222,
    65217,65212,65207,65202,65197,65192,65187,65182,
    65177,65171,65166,65161,65155,65150,65144,65139,
    65133,65128,65122,65117,65111,65105,65099,65094,
    65088,65082,65076,65070,65064,65058,65052,65046,
    65040,65033,65027,65021,65015,65008,65002,64995,
    64989,64982,64976,64969,64963,64956,64949,64943,
    64936,64929,64922,64915,64908,64902,64895,64887,
    64880,64873,64866,64859,64852,64844,64837,64830,
    64822,64815,64808,64800,64793,64785,64777,64770,
    64762,64754,64747,64739,64731,64723,64715,64707,
    64699,64691,64683,64675,64667,64659,64651,64642,
    64634,64626,64617,64609,64600,64592,64584,64575,
    64566,64558,64549,64540,64532,64523,64514,64505,
    64496,64487,64478,64469,64460,64451,64442,64433,
    64424,64414,64405,64396,64387,64377,64368,64358,
    64349,64339,64330,64320,64310,64301,64291,64281,
    64271,64261,64252,64242,64232,64222,64212,64202,
    64192,64181,64171,64161,64151,64140,64130,64120,
    64109,64099,64088,64078,64067,64057,64046,64035,
    64025,64014,64003,63992,63981,63971,63960,63949,
    63938,63927,63915,63904,63893,63882,63871,63859,
    63848,63837,63825,63814,63803,63791,63779,63768,
    63756,63745,63733,63721,63709,63698,63686,63674,
    63662,63650,63638,63626,63614,63602,63590,63578,
    63565,63553,63541,63528,63516,63504,63491,63479,
    63466,63454,63441,63429,63416,63403,63390,63378,
    63365,63352,63339,63326,63313,63300,63287,63274,
    63261,63248,63235,63221,63208,63195,63182,63168,
    63155,63141,63128,63114,63101,63087,63074,63060,
    63046,63032,63019,63005,62991,62977,62963,62949,
    62935,62921,62907,62893,62879,62865,62850,62836,
    62822,62808,62793,62779,62764,62750,62735,62721,
    62706,62692,62677,62662,62648,62633,62618,62603,
    62588,62573,62558,62543,62528,62513,62498,62483,
    62468,62453,62437,62422,62407,62391,62376,62360,
    62345,62329,62314,62298,62283,62267,62251,62236,
    62220,62204,62188,62172,62156,62141,62125,62108,
    62092,62076,62060,62044,62028,62012,61995,61979,
    61963,61946,61930,61913,61897,61880,61864,61847,
    61831,61814,61797,61780,61764,61747,61730,61713,
    61696,61679,61662,61645,61628,61611,61594,61577,
    61559,61542,61525,61507,61490,61473,61455,61438,
    61420,61403,61385,61367,61350,61332,61314,61297,
    61279,61261,61243,61225,61207,61189,61171,61153,
    61135,61117,61099,61081,61062,61044,61026,61007,
    60989,60971,60952,60934,60915,60897,60878,60859,
    60841,60822,60803,60785,60766,60747,60728,60709,
    60690,60671,60652,60633,60614,60595,60576,60556,
    60537,60518,60499,60479,60460,60441,60421,60402,
    60382,60363,60343,60323,60304,60284,60264,60244,
    60225,60205,60185,60165,60145,60125,60105,60085,
    60065,60045,60025,60004,59984,59964,59944,59923,
    59903,59883,59862,59842,59821,59801,59780,59759,
    59739,59718,59697,59677,59656,59635,59614,59593,
    59572,59551,59530,59509,59488,59467,59446,59425,
    59404,59382,59361,59340,59318,59297,59276,59254,
    59233,59211,59190,59168,59146,59125,59103,59081,
    59059,59038,59016,58994,58972,58950,58928,58906,
    58884,58862,58840,58818,58795,58773,58751,58729,
    58706,58684,58662,58639,58617,58594,58572,58549,
    58527,58504,58481,58459,58436,58413,58390,58367,
    58345,58322,58299,58276,58253,58230,58207,58183,
    58160,58137,58114,58091,58067,58044,58021,57997,
    57974,57950,57927,57903,57880,57856,57833,57809,
    57785,57762,57738,57714,57690,57666,57642,57618,
    57594,57570,57546,57522,57498,57474,57450,57426,
    57402,57377,57353,57329,57304,57280,57255,57231,
    57206,57182,57157,57133,57108,57083,57059,57034,
    57009,56984,56959,56935,56910,56885,56860,56835,
    56810,56785,56760,56734,56709,56684,56659,56633,
    56608,56583,56557,56532,56507,56481,56456,56430,
    56404,56379,56353,56328,56302,56276,56250,56225,
    56199,56173,56147,56121,56095,56069,56043,56017,
    55991,55965,55938,55912,55886,55860,55833,55807,
    55781,55754,55728,55701,55675,55648,55622,55595,
    55569,55542,55515,55489,55462,55435,55408,55381,
    55354,55327,55300,55274,55246,55219,55192,55165,
    55138,55111,55084,55056,55029,55002,54974,54947,
    54920,54892,54865,54837,54810,54782,54755,54727,
    54699,54672,54644,54616,54588,54560,54533,54505,
    54477,54449,54421,54393,54365,54337,54308,54280,
    54252,54224,54196,54167,54139,54111,54082,54054,
    54026,53997,53969,53940,53911,53883,53854,53826,
    53797,53768,53739,53711,53682,53653,53624,53595,
    53566,53537,53508,53479,53450,53421,53392,53363,
    53334,53304,53275,53246,53216,53187,53158,53128,
    53099,53069,53040,53010,52981,52951,52922,52892,
    52862,52832,52803,52773,52743,52713,52683,52653,
    52624,52594,52564,52534,52503,52473,52443,52413,
    52383,52353,52322,52292,52262,52231,52201,52171,
    52140,52110,52079,52049,52018,51988,51957,51926,
    51896,51865,51834,51803,51773,51742,51711,51680,
    51649,51618,51587,51556,51525,51494,51463,51432,
    51401,51369,51338,51307,51276,51244,51213,51182,
    51150,51119,51087,51056,51024,50993,50961,50929,
    50898,50866,50834,50803,50771,50739,50707,50675,
    50644,50612,50580,50548,50516,50484,50452,50420,
    50387,50355,50323,50291,50259,50226,50194,50162,
    50129,50097,50065,50032,50000,49967,49935,49902,
    49869,49837,49804,49771,49739,49706,49673,49640,
    49608,49575,49542,49509,49476,49443,49410,49377,
    49344,49311,49278,49244,49211,49178,49145,49112,
    49078,49045,49012,48978,48945,48911,48878,48844,
    48811,48777,48744,48710,48676,48643,48609,48575,
    48542,48508,48474,48440,48406,48372,48338,48304,
    48271,48237,48202,48168,48134,48100,48066,48032,
    47998,47963,47929,47895,47860,47826,47792,47757,
    47723,47688,47654,47619,47585,47550,47516,47481,
    47446,47412,47377,47342,47308,47273,47238,47203,
    47168,47133,47098,47063,47028,46993,46958,46923,
    46888,46853,46818,46783,46747,46712,46677,46642,
    46606,46571,46536,46500,46465,46429,46394,46358,
    46323,46287,46252,46216,46180,46145,46109,46073,
    46037,46002,45966,45930,45894,45858,45822,45786,
    45750,45714,45678,45642,45606,45570,45534,45498,
    45462,45425,45389,45353,45316,45280,45244,45207,
    45171,45135,45098,45062,45025,44989,44952,44915,
    44879,44842,44806,44769,44732,44695,44659,44622,
    44585,44548,44511,44474,44437,44400,44363,44326,
    44289,44252,44215,44178,44141,44104,44067,44029,
    43992,43955,43918,43880,43843,43806,43768,43731,
    43693,43656,43618,43581,43543,43506,43468,43430,
    43393,43355,43317,43280,43242,43204,43166,43128,
    43091,43053,43015,42977,42939,42901,42863,42825,
    42787,42749,42711,42672,42634,42596,42558,42520,
    42481,42443,42405,42366,42328,42290,42251,42213,
    42174,42136,42097,42059,42020,41982,41943,41904,
    41866,41827,41788,41750,41711,41672,41633,41595,
    41556,41517,41478,41439,41400,41361,41322,41283,
    41244,41205,41166,41127,41088,41048,41009,40970,
    40931,40891,40852,40813,40773,40734,40695,40655,
    40616,40576,40537,40497,40458,40418,40379,40339,
    40300,40260,40220,40180,40141,40101,40061,40021,
    39982,39942,39902,39862,39822,39782,39742,39702,
    39662,39622,39582,39542,39502,39462,39422,39382,
    39341,39301,39261,39221,39180,39140,39100,39059,
    39019,38979,38938,38898,38857,38817,38776,38736,
    38695,38655,38614,38573,38533,38492,38451,38411,
    38370,38329,38288,38248,38207,38166,38125,38084,
    38043,38002,37961,37920,37879,37838,37797,37756,
    37715,37674,37633,37592,37551,37509,37468,37427,
    37386,37344,37303,37262,37220,37179,37137,37096,
    37055,37013,36972,36930,36889,36847,36805,36764,
    36722,36681,36639,36597,36556,36514,36472,36430,
    36388,36347,36305,36263,36221,36179,36137,36095,
    36053,36011,35969,35927,35885,35843,35801,35759,
    35717,35675,35633,35590,35548,35506,35464,35421,
    35379,35337,35294,35252,35210,35167,35125,35082,
    35040,34997,34955,34912,34870,34827,34785,34742,
    34699,34657,34614,34571,34529,34486,34443,34400,
    34358,34315,34272,34229,34186,34143,34100,34057,
    34015,33972,33929,33886,33843,33799,33756,33713,
    33670,33627,33584,33541,33498,33454,33411,33368,
    33325,33281,33238,33195,33151,33108,33065,33021,
    32978,32934,32891,32847,32804,32760,32717,32673,
    32630,32586,32542,32499,32455,32411,32368,32324,
    32280,32236,32193,32149,32105,32061,32017,31974,
    31930,31886,31842,31798,31754,31710,31666,31622,
    31578,31534,31490,31446,31402,31357,31313,31269,
    31225,31181,31136,31092,31048,31004,30959,30915,
    30871,30826,30782,30738,30693,30649,30604,30560,
    30515,30471,30426,30382,30337,30293,30248,30204,
    30159,30114,30070,30025,29980,29936,29891,29846,
    29801,29757,29712,29667,29622,29577,29533,29488,
    29443,29398,29353,29308,29263,29218,29173,29128,
    29083,29038,28993,28948,28903,28858,28812,28767,
    28722,28677,28632,28586,28541,28496,28451,28405,
    28360,28315,28269,28224,28179,28133,28088,28042,
    27997,27952,27906,27861,27815,27770,27724,27678,
    27633,27587,27542,27496,27450,27405,27359,27313,
    27268,27222,27176,27131,27085,27039,26993,26947,
    26902,26856,26810,26764,26718,26672,26626,26580,
    26534,26488,26442,26396,26350,26304,26258,26212,
    26166,26120,26074,26028,25982,25936,25889,25843,
    25797,25751,25705,25658,25612,25566,25520,25473,
    25427,25381,25334,25288,25241,25195,25149,25102,
    25056,25009,24963,24916,24870,24823,24777,24730,
    24684,24637,24591,24544,24497,24451,24404,24357,
    24311,24264,24217,24171,24124,24077,24030,23984,
    23937,23890,23843,23796,23750,23703,23656,23609,
    23562,23515,23468,23421,23374,23327,23280,23233,
    23186,23139,23092,23045,22998,22951,22904,22857,
    22810,22763,22716,22668,22621,22574,22527,22480,
    22433,22385,22338,22291,22243,22196,22149,22102,
    22054,22007,21960,21912,21865,21817,21770,21723,
    21675,21628,21580,21533,21485,21438,21390,21343,
    21295,21248,21200,21153,21105,21057,21010,20962,
    20915,20867,20819,20772,20724,20676,20629,20581,
    20533,20485,20438,20390,20342,20294,20246,20199,
    20151,20103,20055,20007,19959,19912,19864,19816,
    19768,19720,19672,19624,19576,19528,19480,19432,
    19384,19336,19288,19240,19192,19144,19096,19048,
    19000,18951,18903,18855,18807,18759,18711,18663,
    18614,18566,18518,18470,18421,18373,18325,18277,
    18228,18180,18132,18084,18035,17987,17939,17890,
    17842,17793,17745,17697,17648,17600,17551,17503,
    17455,17406,17358,17309,17261,17212,17164,17115,
    17067,17018,16970,16921,16872,16824,16775,16727,
    16678,16629,16581,16532,16484,16435,16386,16338,
    16289,16240,16191,16143,16094,16045,15997,15948,
    15899,15850,15802,15753,15704,15655,15606,15557,
    15509,15460,15411,15362,15313,15264,15215,15167,
    15118,15069,15020,14971,14922,14873,14824,14775,
    14726,14677,14628,14579,14530,14481,14432,14383,
    14334,14285,14236,14187,14138,14089,14040,13990,
    13941,13892,13843,13794,13745,13696,13646,13597,
    13548,13499,13450,13401,13351,13302,13253,13204,
    13154,13105,13056,13007,12957,12908,12859,12810,
    12760,12711,12662,12612,12563,12514,12464,12415,
    12366,12316,12267,12218,12168,12119,12069,12020,
    11970,11921,11872,11822,11773,11723,11674,11624,
    11575,11525,11476,11426,11377,11327,11278,11228,
    11179,11129,11080,11030,10981,10931,10882,10832,
    10782,10733,10683,10634,10584,10534,10485,10435,
    10386,10336,10286,10237,10187,10137,10088,10038,
    9988,9939,9889,9839,9790,9740,9690,9640,
    9591,9541,9491,9442,9392,9342,9292,9243,
    9193,9143,9093,9043,8994,8944,8894,8844,
    8794,8745,8695,8645,8595,8545,8496,8446,
    8396,8346,8296,8246,8196,8147,8097,8047,
    7997,7947,7897,7847,7797,7747,7697,7648,
    7598,7548,7498,7448,7398,7348,7298,7248,
    7198,7148,7098,7048,6998,6948,6898,6848,
    6798,6748,6698,6648,6598,6548,6498,6448,
    6398,6348,6298,6248,6198,6148,6098,6048,
    5998,5948,5898,5848,5798,5748,5697,5647,
    5597,5547,5497,5447,5397,5347,5297,5247,
    5197,5146,5096,5046,4996,4946,4896,4846,
    4796,4745,4695,4645,4595,4545,4495,4445,
    4394,4344,4294,4244,4194,4144,4093,4043,
    3993,3943,3893,3843,3792,3742,3692,3642,
    3592,3541,3491,3441,3391,3341,3291,3240,
    3190,3140,3090,3039,2989,2939,2889,2839,
    2788,2738,2688,2638,2587,2537,2487,2437,
    2387,2336,2286,2236,2186,2135,2085,2035,
    1985,1934,1884,1834,1784,1733,1683,1633,
    1583,1532,1482,1432,1382,1331,1281,1231,
    1181,1130,1080,1030,980,929,879,829,
    779,728,678,628,578,527,477,427,
    376,326,276,226,175,125,75,25,
    -25,-75,-125,-175,-226,-276,-326,-376,
    -427,-477,-527,-578,-628,-678,-728,-779,
    -829,-879,-929,-980,-1030,-1080,-1130,-1181,
    -1231,-1281,-1331,-1382,-1432,-1482,-1532,-1583,
    -1633,-1683,-1733,-1784,-1834,-1884,-1934,-1985,
    -2035,-2085,-2135,-2186,-2236,-2286,-2336,-2387,
    -2437,-2487,-2537,-2588,-2638,-2688,-2738,-2788,
    -2839,-2889,-2939,-2989,-3039,-3090,-3140,-3190,
    -3240,-3291,-3341,-3391,-3441,-3491,-3541,-3592,
    -3642,-3692,-3742,-3792,-3843,-3893,-3943,-3993,
    -4043,-4093,-4144,-4194,-4244,-4294,-4344,-4394,
    -4445,-4495,-4545,-4595,-4645,-4695,-4745,-4796,
    -4846,-4896,-4946,-4996,-5046,-5096,-5146,-5197,
    -5247,-5297,-5347,-5397,-5447,-5497,-5547,-5597,
    -5647,-5697,-5748,-5798,-5848,-5898,-5948,-5998,
    -6048,-6098,-6148,-6198,-6248,-6298,-6348,-6398,
    -6448,-6498,-6548,-6598,-6648,-6698,-6748,-6798,
    -6848,-6898,-6948,-6998,-7048,-7098,-7148,-7198,
    -7248,-7298,-7348,-7398,-7448,-7498,-7548,-7598,
    -7648,-7697,-7747,-7797,-7847,-7897,-7947,-7997,
    -8047,-8097,-8147,-8196,-8246,-8296,-8346,-8396,
    -8446,-8496,-8545,-8595,-8645,-8695,-8745,-8794,
    -8844,-8894,-8944,-8994,-9043,-9093,-9143,-9193,
    -9243,-9292,-9342,-9392,-9442,-9491,-9541,-9591,
    -9640,-9690,-9740,-9790,-9839,-9889,-9939,-9988,
    -10038,-10088,-10137,-10187,-10237,-10286,-10336,-10386,
    -10435,-10485,-10534,-10584,-10634,-10683,-10733,-10782,
    -10832,-10882,-10931,-10981,-11030,-11080,-11129,-11179,
    -11228,-11278,-11327,-11377,-11426,-11476,-11525,-11575,
    -11624,-11674,-11723,-11773,-11822,-11872,-11921,-11970,
    -12020,-12069,-12119,-12168,-12218,-12267,-12316,-12366,
    -12415,-12464,-12514,-12563,-12612,-12662,-12711,-12760,
    -12810,-12859,-12908,-12957,-13007,-13056,-13105,-13154,
    -13204,-13253,-13302,-13351,-13401,-13450,-13499,-13548,
    -13597,-13647,-13696,-13745,-13794,-13843,-13892,-13941,
    -13990,-14040,-14089,-14138,-14187,-14236,-14285,-14334,
    -14383,-14432,-14481,-14530,-14579,-14628,-14677,-14726,
    -14775,-14824,-14873,-14922,-14971,-15020,-15069,-15118,
    -15167,-15215,-15264,-15313,-15362,-15411,-15460,-15509,
    -15557,-15606,-15655,-15704,-15753,-15802,-15850,-15899,
    -15948,-15997,-16045,-16094,-16143,-16191,-16240,-16289,
    -16338,-16386,-16435,-16484,-16532,-16581,-16629,-16678,
    -16727,-16775,-16824,-16872,-16921,-16970,-17018,-17067,
    -17115,-17164,-17212,-17261,-17309,-17358,-17406,-17455,
    -17503,-17551,-17600,-17648,-17697,-17745,-17793,-17842,
    -17890,-17939,-17987,-18035,-18084,-18132,-18180,-18228,
    -18277,-18325,-18373,-18421,-18470,-18518,-18566,-18614,
    -18663,-18711,-18759,-18807,-18855,-18903,-18951,-19000,
    -19048,-19096,-19144,-19192,-19240,-19288,-19336,-19384,
    -19432,-19480,-19528,-19576,-19624,-19672,-19720,-19768,
    -19816,-19864,-19912,-19959,-20007,-20055,-20103,-20151,
    -20199,-20246,-20294,-20342,-20390,-20438,-20485,-20533,
    -20581,-20629,-20676,-20724,-20772,-20819,-20867,-20915,
    -20962,-21010,-21057,-21105,-21153,-21200,-21248,-21295,
    -21343,-21390,-21438,-21485,-21533,-21580,-21628,-21675,
    -21723,-21770,-21817,-21865,-21912,-21960,-22007,-22054,
    -22102,-22149,-22196,-22243,-22291,-22338,-22385,-22433,
    -22480,-22527,-22574,-22621,-22668,-22716,-22763,-22810,
    -22857,-22904,-22951,-22998,-23045,-23092,-23139,-23186,
    -23233,-23280,-23327,-23374,-23421,-23468,-23515,-23562,
    -23609,-23656,-23703,-23750,-23796,-23843,-23890,-23937,
    -23984,-24030,-24077,-24124,-24171,-24217,-24264,-24311,
    -24357,-24404,-24451,-24497,-24544,-24591,-24637,-24684,
    -24730,-24777,-24823,-24870,-24916,-24963,-25009,-25056,
    -25102,-25149,-25195,-25241,-25288,-25334,-25381,-25427,
    -25473,-25520,-25566,-25612,-25658,-25705,-25751,-25797,
    -25843,-25889,-25936,-25982,-26028,-26074,-26120,-26166,
    -26212,-26258,-26304,-26350,-26396,-26442,-26488,-26534,
    -26580,-26626,-26672,-26718,-26764,-26810,-26856,-26902,
    -26947,-26993,-27039,-27085,-27131,-27176,-27222,-27268,
    -27313,-27359,-27405,-27450,-27496,-27542,-27587,-27633,
    -27678,-27724,-27770,-27815,-27861,-27906,-27952,-27997,
    -28042,-28088,-28133,-28179,-28224,-28269,-28315,-28360,
    -28405,-28451,-28496,-28541,-28586,-28632,-28677,-28722,
    -28767,-28812,-28858,-28903,-28948,-28993,-29038,-29083,
    -29128,-29173,-29218,-29263,-29308,-29353,-29398,-29443,
    -29488,-29533,-29577,-29622,-29667,-29712,-29757,-29801,
    -29846,-29891,-29936,-29980,-30025,-30070,-30114,-30159,
    -30204,-30248,-30293,-30337,-30382,-30426,-30471,-30515,
    -30560,-30604,-30649,-30693,-30738,-30782,-30826,-30871,
    -30915,-30959,-31004,-31048,-31092,-31136,-31181,-31225,
    -31269,-31313,-31357,-31402,-31446,-31490,-31534,-31578,
    -31622,-31666,-31710,-31754,-31798,-31842,-31886,-31930,
    -31974,-32017,-32061,-32105,-32149,-32193,-32236,-32280,
    -32324,-32368,-32411,-32455,-32499,-32542,-32586,-32630,
    -32673,-32717,-32760,-32804,-32847,-32891,-32934,-32978,
    -33021,-33065,-33108,-33151,-33195,-33238,-33281,-33325,
    -33368,-33411,-33454,-33498,-33541,-33584,-33627,-33670,
    -33713,-33756,-33799,-33843,-33886,-33929,-33972,-34015,
    -34057,-34100,-34143,-34186,-34229,-34272,-34315,-34358,
    -34400,-34443,-34486,-34529,-34571,-34614,-34657,-34699,
    -34742,-34785,-34827,-34870,-34912,-34955,-34997,-35040,
    -35082,-35125,-35167,-35210,-35252,-35294,-35337,-35379,
    -35421,-35464,-35506,-35548,-35590,-35633,-35675,-35717,
    -35759,-35801,-35843,-35885,-35927,-35969,-36011,-36053,
    -36095,-36137,-36179,-36221,-36263,-36305,-36347,-36388,
    -36430,-36472,-36514,-36555,-36597,-36639,-36681,-36722,
    -36764,-36805,-36847,-36889,-36930,-36972,-37013,-37055,
    -37096,-37137,-37179,-37220,-37262,-37303,-37344,-37386,
    -37427,-37468,-37509,-37551,-37592,-37633,-37674,-37715,
    -37756,-37797,-37838,-37879,-37920,-37961,-38002,-38043,
    -38084,-38125,-38166,-38207,-38248,-38288,-38329,-38370,
    -38411,-38451,-38492,-38533,-38573,-38614,-38655,-38695,
    -38736,-38776,-38817,-38857,-38898,-38938,-38979,-39019,
    -39059,-39100,-39140,-39180,-39221,-39261,-39301,-39341,
    -39382,-39422,-39462,-39502,-39542,-39582,-39622,-39662,
    -39702,-39742,-39782,-39822,-39862,-39902,-39942,-39982,
    -40021,-40061,-40101,-40141,-40180,-40220,-40260,-40299,
    -40339,-40379,-40418,-40458,-40497,-40537,-40576,-40616,
    -40655,-40695,-40734,-40773,-40813,-40852,-40891,-40931,
    -40970,-41009,-41048,-41087,-41127,-41166,-41205,-41244,
    -41283,-41322,-41361,-41400,-41439,-41478,-41517,-41556,
    -41595,-41633,-41672,-41711,-41750,-41788,-41827,-41866,
    -41904,-41943,-41982,-42020,-42059,-42097,-42136,-42174,
    -42213,-42251,-42290,-42328,-42366,-42405,-42443,-42481,
    -42520,-42558,-42596,-42634,-42672,-42711,-42749,-42787,
    -42825,-42863,-42901,-42939,-42977,-43015,-43053,-43091,
    -43128,-43166,-43204,-43242,-43280,-43317,-43355,-43393,
    -43430,-43468,-43506,-43543,-43581,-43618,-43656,-43693,
    -43731,-43768,-43806,-43843,-43880,-43918,-43955,-43992,
    -44029,-44067,-44104,-44141,-44178,-44215,-44252,-44289,
    -44326,-44363,-44400,-44437,-44474,-44511,-44548,-44585,
    -44622,-44659,-44695,-44732,-44769,-44806,-44842,-44879,
    -44915,-44952,-44989,-45025,-45062,-45098,-45135,-45171,
    -45207,-45244,-45280,-45316,-45353,-45389,-45425,-45462,
    -45498,-45534,-45570,-45606,-45642,-45678,-45714,-45750,
    -45786,-45822,-45858,-45894,-45930,-45966,-46002,-46037,
    -46073,-46109,-46145,-46180,-46216,-46252,-46287,-46323,
    -46358,-46394,-46429,-46465,-46500,-46536,-46571,-46606,
    -46642,-46677,-46712,-46747,-46783,-46818,-46853,-46888,
    -46923,-46958,-46993,-47028,-47063,-47098,-47133,-47168,
    -47203,-47238,-47273,-47308,-47342,-47377,-47412,-47446,
    -47481,-47516,-47550,-47585,-47619,-47654,-47688,-47723,
    -47757,-47792,-47826,-47860,-47895,-47929,-47963,-47998,
    -48032,-48066,-48100,-48134,-48168,-48202,-48236,-48271,
    -48304,-48338,-48372,-48406,-48440,-48474,-48508,-48542,
    -48575,-48609,-48643,-48676,-48710,-48744,-48777,-48811,
    -48844,-48878,-48911,-48945,-48978,-49012,-49045,-49078,
    -49112,-49145,-49178,-49211,-49244,-49278,-49311,-49344,
    -49377,-49410,-49443,-49476,-49509,-49542,-49575,-49608,
    -49640,-49673,-49706,-49739,-49771,-49804,-49837,-49869,
    -49902,-49935,-49967,-50000,-50032,-50065,-50097,-50129,
    -50162,-50194,-50226,-50259,-50291,-50323,-50355,-50387,
    -50420,-50452,-50484,-50516,-50548,-50580,-50612,-50644,
    -50675,-50707,-50739,-50771,-50803,-50834,-50866,-50898,
    -50929,-50961,-50993,-51024,-51056,-51087,-51119,-51150,
    -51182,-51213,-51244,-51276,-51307,-51338,-51369,-51401,
    -51432,-51463,-51494,-51525,-51556,-51587,-51618,-51649,
    -51680,-51711,-51742,-51773,-51803,-51834,-51865,-51896,
    -51926,-51957,-51988,-52018,-52049,-52079,-52110,-52140,
    -52171,-52201,-52231,-52262,-52292,-52322,-52353,-52383,
    -52413,-52443,-52473,-52503,-52534,-52564,-52594,-52624,
    -52653,-52683,-52713,-52743,-52773,-52803,-52832,-52862,
    -52892,-52922,-52951,-52981,-53010,-53040,-53069,-53099,
    -53128,-53158,-53187,-53216,-53246,-53275,-53304,-53334,
    -53363,-53392,-53421,-53450,-53479,-53508,-53537,-53566,
    -53595,-53624,-53653,-53682,-53711,-53739,-53768,-53797,
    -53826,-53854,-53883,-53911,-53940,-53969,-53997,-54026,
    -54054,-54082,-54111,-54139,-54167,-54196,-54224,-54252,
    -54280,-54308,-54337,-54365,-54393,-54421,-54449,-54477,
    -54505,-54533,-54560,-54588,-54616,-54644,-54672,-54699,
    -54727,-54755,-54782,-54810,-54837,-54865,-54892,-54920,
    -54947,-54974,-55002,-55029,-55056,-55084,-55111,-55138,
    -55165,-55192,-55219,-55246,-55274,-55300,-55327,-55354,
    -55381,-55408,-55435,-55462,-55489,-55515,-55542,-55569,
    -55595,-55622,-55648,-55675,-55701,-55728,-55754,-55781,
    -55807,-55833,-55860,-55886,-55912,-55938,-55965,-55991,
    -56017,-56043,-56069,-56095,-56121,-56147,-56173,-56199,
    -56225,-56250,-56276,-56302,-56328,-56353,-56379,-56404,
    -56430,-56456,-56481,-56507,-56532,-56557,-56583,-56608,
    -56633,-56659,-56684,-56709,-56734,-56760,-56785,-56810,
    -56835,-56860,-56885,-56910,-56935,-56959,-56984,-57009,
    -57034,-57059,-57083,-57108,-57133,-57157,-57182,-57206,
    -57231,-57255,-57280,-57304,-57329,-57353,-57377,-57402,
    -57426,-57450,-57474,-57498,-57522,-57546,-57570,-57594,
    -57618,-57642,-57666,-57690,-57714,-57738,-57762,-57785,
    -57809,-57833,-57856,-57880,-57903,-57927,-57950,-57974,
    -57997,-58021,-58044,-58067,-58091,-58114,-58137,-58160,
    -58183,-58207,-58230,-58253,-58276,-58299,-58322,-58345,
    -58367,-58390,-58413,-58436,-58459,-58481,-58504,-58527,
    -58549,-58572,-58594,-58617,-58639,-58662,-58684,-58706,
    -58729,-58751,-58773,-58795,-58818,-58840,-58862,-58884,
    -58906,-58928,-58950,-58972,-58994,-59016,-59038,-59059,
    -59081,-59103,-59125,-59146,-59168,-59190,-59211,-59233,
    -59254,-59276,-59297,-59318,-59340,-59361,-59382,-59404,
    -59425,-59446,-59467,-59488,-59509,-59530,-59551,-59572,
    -59593,-59614,-59635,-59656,-59677,-59697,-59718,-59739,
    -59759,-59780,-59801,-59821,-59842,-59862,-59883,-59903,
    -59923,-59944,-59964,-59984,-60004,-60025,-60045,-60065,
    -60085,-60105,-60125,-60145,-60165,-60185,-60205,-60225,
    -60244,-60264,-60284,-60304,-60323,-60343,-60363,-60382,
    -60402,-60421,-60441,-60460,-60479,-60499,-60518,-60537,
    -60556,-60576,-60595,-60614,-60633,-60652,-60671,-60690,
    -60709,-60728,-60747,-60766,-60785,-60803,-60822,-60841,
    -60859,-60878,-60897,-60915,-60934,-60952,-60971,-60989,
    -61007,-61026,-61044,-61062,-61081,-61099,-61117,-61135,
    -61153,-61171,-61189,-61207,-61225,-61243,-61261,-61279,
    -61297,-61314,-61332,-61350,-61367,-61385,-61403,-61420,
    -61438,-61455,-61473,-61490,-61507,-61525,-61542,-61559,
    -61577,-61594,-61611,-61628,-61645,-61662,-61679,-61696,
    -61713,-61730,-61747,-61764,-61780,-61797,-61814,-61831,
    -61847,-61864,-61880,-61897,-61913,-61930,-61946,-61963,
    -61979,-61995,-62012,-62028,-62044,-62060,-62076,-62092,
    -62108,-62125,-62141,-62156,-62172,-62188,-62204,-62220,
    -62236,-62251,-62267,-62283,-62298,-62314,-62329,-62345,
    -62360,-62376,-62391,-62407,-62422,-62437,-62453,-62468,
    -62483,-62498,-62513,-62528,-62543,-62558,-62573,-62588,
    -62603,-62618,-62633,-62648,-62662,-62677,-62692,-62706,
    -62721,-62735,-62750,-62764,-62779,-62793,-62808,-62822,
    -62836,-62850,-62865,-62879,-62893,-62907,-62921,-62935,
    -62949,-62963,-62977,-62991,-63005,-63019,-63032,-63046,
    -63060,-63074,-63087,-63101,-63114,-63128,-63141,-63155,
    -63168,-63182,-63195,-63208,-63221,-63235,-63248,-63261,
    -63274,-63287,-63300,-63313,-63326,-63339,-63352,-63365,
    -63378,-63390,-63403,-63416,-63429,-63441,-63454,-63466,
    -63479,-63491,-63504,-63516,-63528,-63541,-63553,-63565,
    -63578,-63590,-63602,-63614,-63626,-63638,-63650,-63662,
    -63674,-63686,-63698,-63709,-63721,-63733,-63745,-63756,
    -63768,-63779,-63791,-63803,-63814,-63825,-63837,-63848,
    -63859,-63871,-63882,-63893,-63904,-63915,-63927,-63938,
    -63949,-63960,-63971,-63981,-63992,-64003,-64014,-64025,
    -64035,-64046,-64057,-64067,-64078,-64088,-64099,-64109,
    -64120,-64130,-64140,-64151,-64161,-64171,-64181,-64192,
    -64202,-64212,-64222,-64232,-64242,-64252,-64261,-64271,
    -64281,-64291,-64301,-64310,-64320,-64330,-64339,-64349,
    -64358,-64368,-64377,-64387,-64396,-64405,-64414,-64424,
    -64433,-64442,-64451,-64460,-64469,-64478,-64487,-64496,
    -64505,-64514,-64523,-64532,-64540,-64549,-64558,-64566,
    -64575,-64584,-64592,-64601,-64609,-64617,-64626,-64634,
    -64642,-64651,-64659,-64667,-64675,-64683,-64691,-64699,
    -64707,-64715,-64723,-64731,-64739,-64747,-64754,-64762,
    -64770,-64777,-64785,-64793,-64800,-64808,-64815,-64822,
    -64830,-64837,-64844,-64852,-64859,-64866,-64873,-64880,
    -64887,-64895,-64902,-64908,-64915,-64922,-64929,-64936,
    -64943,-64949,-64956,-64963,-64969,-64976,-64982,-64989,
    -64995,-65002,-65008,-65015,-65021,-65027,-65033,-65040,
    -65046,-65052,-65058,-65064,-65070,-65076,-65082,-65088,
    -65094,-65099,-65105,-65111,-65117,-65122,-65128,-65133,
    -65139,-65144,-65150,-65155,-65161,-65166,-65171,-65177,
    -65182,-65187,-65192,-65197,-65202,-65207,-65212,-65217,
    -65222,-65227,-65232,-65237,-65242,-65246,-65251,-65256,
    -65260,-65265,-65270,-65274,-65279,-65283,-65287,-65292,
    -65296,-65300,-65305,-65309,-65313,-65317,-65321,-65325,
    -65329,-65333,-65337,-65341,-65345,-65349,-65352,-65356,
    -65360,-65363,-65367,-65371,-65374,-65378,-65381,-65385,
    -65388,-65391,-65395,-65398,-65401,-65404,-65408,-65411,
    -65414,-65417,-65420,-65423,-65426,-65429,-65431,-65434,
    -65437,-65440,-65442,-65445,-65448,-65450,-65453,-65455,
    -65458,-65460,-65463,-65465,-65467,-65470,-65472,-65474,
    -65476,-65478,-65480,-65482,-65484,-65486,-65488,-65490,
    -65492,-65494,-65496,-65497,-65499,-65501,-65502,-65504,
    -65505,-65507,-65508,-65510,-65511,-65513,-65514,-65515,
    -65516,-65518,-65519,-65520,-65521,-65522,-65523,-65524,
    -65525,-65526,-65527,-65527,-65528,-65529,-65530,-65530,
    -65531,-65531,-65532,-65532,-65533,-65533,-65534,-65534,
    -65534,-65535,-65535,-65535,-65535,-65535,-65535,-65535,
    -65535,-65535,-65535,-65535,-65535,-65535,-65535,-65534,
    -65534,-65534,-65533,-65533,-65532,-65532,-65531,-65531,
    -65530,-65530,-65529,-65528,-65527,-65527,-65526,-65525,
    -65524,-65523,-65522,-65521,-65520,-65519,-65518,-65516,
    -65515,-65514,-65513,-65511,-65510,-65508,-65507,-65505,
    -65504,-65502,-65501,-65499,-65497,-65496,-65494,-65492,
    -65490,-65488,-65486,-65484,-65482,-65480,-65478,-65476,
    -65474,-65472,-65470,-65467,-65465,-65463,-65460,-65458,
    -65455,-65453,-65450,-65448,-65445,-65442,-65440,-65437,
    -65434,-65431,-65429,-65426,-65423,-65420,-65417,-65414,
    -65411,-65408,-65404,-65401,-65398,-65395,-65391,-65388,
    -65385,-65381,-65378,-65374,-65371,-65367,-65363,-65360,
    -65356,-65352,-65349,-65345,-65341,-65337,-65333,-65329,
    -65325,-65321,-65317,-65313,-65309,-65305,-65300,-65296,
    -65292,-65287,-65283,-65279,-65274,-65270,-65265,-65260,
    -65256,-65251,-65246,-65242,-65237,-65232,-65227,-65222,
    -65217,-65212,-65207,-65202,-65197,-65192,-65187,-65182,
    -65177,-65171,-65166,-65161,-65155,-65150,-65144,-65139,
    -65133,-65128,-65122,-65117,-65111,-65105,-65099,-65094,
    -65088,-65082,-65076,-65070,-65064,-65058,-65052,-65046,
    -65040,-65033,-65027,-65021,-65015,-65008,-65002,-64995,
    -64989,-64982,-64976,-64969,-64963,-64956,-64949,-64943,
    -64936,-64929,-64922,-64915,-64908,-64902,-64895,-64887,
    -64880,-64873,-64866,-64859,-64852,-64844,-64837,-64830,
    -64822,-64815,-64808,-64800,-64793,-64785,-64777,-64770,
    -64762,-64754,-64747,-64739,-64731,-64723,-64715,-64707,
    -64699,-64691,-64683,-64675,-64667,-64659,-64651,-64642,
    -64634,-64626,-64617,-64609,-64601,-64592,-64584,-64575,
    -64566,-64558,-64549,-64540,-64532,-64523,-64514,-64505,
    -64496,-64487,-64478,-64469,-64460,-64451,-64442,-64433,
    -64424,-64414,-64405,-64396,-64387,-64377,-64368,-64358,
    -64349,-64339,-64330,-64320,-64310,-64301,-64291,-64281,
    -64271,-64261,-64252,-64242,-64232,-64222,-64212,-64202,
    -64192,-64181,-64171,-64161,-64151,-64140,-64130,-64120,
    -64109,-64099,-64088,-64078,-64067,-64057,-64046,-64035,
    -64025,-64014,-64003,-63992,-63981,-63971,-63960,-63949,
    -63938,-63927,-63915,-63904,-63893,-63882,-63871,-63859,
    -63848,-63837,-63825,-63814,-63803,-63791,-63779,-63768,
    -63756,-63745,-63733,-63721,-63709,-63698,-63686,-63674,
    -63662,-63650,-63638,-63626,-63614,-63602,-63590,-63578,
    -63565,-63553,-63541,-63528,-63516,-63504,-63491,-63479,
    -63466,-63454,-63441,-63429,-63416,-63403,-63390,-63378,
    -63365,-63352,-63339,-63326,-63313,-63300,-63287,-63274,
    -63261,-63248,-63235,-63221,-63208,-63195,-63182,-63168,
    -63155,-63141,-63128,-63114,-63101,-63087,-63074,-63060,
    -63046,-63032,-63019,-63005,-62991,-62977,-62963,-62949,
    -62935,-62921,-62907,-62893,-62879,-62865,-62850,-62836,
    -62822,-62808,-62793,-62779,-62764,-62750,-62735,-62721,
    -62706,-62692,-62677,-62662,-62648,-62633,-62618,-62603,
    -62588,-62573,-62558,-62543,-62528,-62513,-62498,-62483,
    -62468,-62453,-62437,-62422,-62407,-62391,-62376,-62360,
    -62345,-62329,-62314,-62298,-62283,-62267,-62251,-62236,
    -62220,-62204,-62188,-62172,-62156,-62141,-62125,-62108,
    -62092,-62076,-62060,-62044,-62028,-62012,-61995,-61979,
    -61963,-61946,-61930,-61913,-61897,-61880,-61864,-61847,
    -61831,-61814,-61797,-61780,-61764,-61747,-61730,-61713,
    -61696,-61679,-61662,-61645,-61628,-61611,-61594,-61577,
    -61559,-61542,-61525,-61507,-61490,-61473,-61455,-61438,
    -61420,-61403,-61385,-61367,-61350,-61332,-61314,-61297,
    -61279,-61261,-61243,-61225,-61207,-61189,-61171,-61153,
    -61135,-61117,-61099,-61081,-61062,-61044,-61026,-61007,
    -60989,-60971,-60952,-60934,-60915,-60897,-60878,-60859,
    -60841,-60822,-60803,-60785,-60766,-60747,-60728,-60709,
    -60690,-60671,-60652,-60633,-60614,-60595,-60576,-60556,
    -60537,-60518,-60499,-60479,-60460,-60441,-60421,-60402,
    -60382,-60363,-60343,-60323,-60304,-60284,-60264,-60244,
    -60225,-60205,-60185,-60165,-60145,-60125,-60105,-60085,
    -60065,-60045,-60025,-60004,-59984,-59964,-59944,-59923,
    -59903,-59883,-59862,-59842,-59821,-59801,-59780,-59759,
    -59739,-59718,-59697,-59677,-59656,-59635,-59614,-59593,
    -59572,-59551,-59530,-59509,-59488,-59467,-59446,-59425,
    -59404,-59382,-59361,-59340,-59318,-59297,-59276,-59254,
    -59233,-59211,-59189,-59168,-59146,-59125,-59103,-59081,
    -59059,-59038,-59016,-58994,-58972,-58950,-58928,-58906,
    -58884,-58862,-58840,-58818,-58795,-58773,-58751,-58729,
    -58706,-58684,-58662,-58639,-58617,-58594,-58572,-58549,
    -58527,-58504,-58481,-58459,-58436,-58413,-58390,-58367,
    -58345,-58322,-58299,-58276,-58253,-58230,-58207,-58183,
    -58160,-58137,-58114,-58091,-58067,-58044,-58021,-57997,
    -57974,-57950,-57927,-57903,-57880,-57856,-57833,-57809,
    -57785,-57762,-57738,-57714,-57690,-57666,-57642,-57618,
    -57594,-57570,-57546,-57522,-57498,-57474,-57450,-57426,
    -57402,-57377,-57353,-57329,-57304,-57280,-57255,-57231,
    -57206,-57182,-57157,-57133,-57108,-57083,-57059,-57034,
    -57009,-56984,-56959,-56935,-56910,-56885,-56860,-56835,
    -56810,-56785,-56760,-56734,-56709,-56684,-56659,-56633,
    -56608,-56583,-56557,-56532,-56507,-56481,-56456,-56430,
    -56404,-56379,-56353,-56328,-56302,-56276,-56250,-56225,
    -56199,-56173,-56147,-56121,-56095,-56069,-56043,-56017,
    -55991,-55965,-55938,-55912,-55886,-55860,-55833,-55807,
    -55781,-55754,-55728,-55701,-55675,-55648,-55622,-55595,
    -55569,-55542,-55515,-55489,-55462,-55435,-55408,-55381,
    -55354,-55327,-55300,-55274,-55246,-55219,-55192,-55165,
    -55138,-55111,-55084,-55056,-55029,-55002,-54974,-54947,
    -54920,-54892,-54865,-54837,-54810,-54782,-54755,-54727,
    -54699,-54672,-54644,-54616,-54588,-54560,-54533,-54505,
    -54477,-54449,-54421,-54393,-54365,-54337,-54308,-54280,
    -54252,-54224,-54196,-54167,-54139,-54111,-54082,-54054,
    -54026,-53997,-53969,-53940,-53911,-53883,-53854,-53826,
    -53797,-53768,-53739,-53711,-53682,-53653,-53624,-53595,
    -53566,-53537,-53508,-53479,-53450,-53421,-53392,-53363,
    -53334,-53304,-53275,-53246,-53216,-53187,-53158,-53128,
    -53099,-53069,-53040,-53010,-52981,-52951,-52922,-52892,
    -52862,-52832,-52803,-52773,-52743,-52713,-52683,-52653,
    -52624,-52594,-52564,-52534,-52503,-52473,-52443,-52413,
    -52383,-52353,-52322,-52292,-52262,-52231,-52201,-52171,
    -52140,-52110,-52079,-52049,-52018,-51988,-51957,-51926,
    -51896,-51865,-51834,-51803,-51773,-51742,-51711,-51680,
    -51649,-51618,-51587,-51556,-51525,-51494,-51463,-51432,
    -51401,-51369,-51338,-51307,-51276,-51244,-51213,-51182,
    -51150,-51119,-51087,-51056,-51024,-50993,-50961,-50929,
    -50898,-50866,-50834,-50803,-50771,-50739,-50707,-50675,
    -50644,-50612,-50580,-50548,-50516,-50484,-50452,-50420,
    -50387,-50355,-50323,-50291,-50259,-50226,-50194,-50162,
    -50129,-50097,-50065,-50032,-50000,-49967,-49935,-49902,
    -49869,-49837,-49804,-49771,-49739,-49706,-49673,-49640,
    -49608,-49575,-49542,-49509,-49476,-49443,-49410,-49377,
    -49344,-49311,-49278,-49244,-49211,-49178,-49145,-49112,
    -49078,-49045,-49012,-48978,-48945,-48911,-48878,-48844,
    -48811,-48777,-48744,-48710,-48676,-48643,-48609,-48575,
    -48542,-48508,-48474,-48440,-48406,-48372,-48338,-48305,
    -48271,-48237,-48202,-48168,-48134,-48100,-48066,-48032,
    -47998,-47963,-47929,-47895,-47860,-47826,-47792,-47757,
    -47723,-47688,-47654,-47619,-47585,-47550,-47516,-47481,
    -47446,-47412,-47377,-47342,-47307,-47273,-47238,-47203,
    -47168,-47133,-47098,-47063,-47028,-46993,-46958,-46923,
    -46888,-46853,-46818,-46783,-46747,-46712,-46677,-46642,
    -46606,-46571,-46536,-46500,-46465,-46429,-46394,-46358,
    -46323,-46287,-46251,-46216,-46180,-46145,-46109,-46073,
    -46037,-46002,-45966,-45930,-45894,-45858,-45822,-45786,
    -45750,-45714,-45678,-45642,-45606,-45570,-45534,-45498,
    -45462,-45425,-45389,-45353,-45316,-45280,-45244,-45207,
    -45171,-45135,-45098,-45062,-45025,-44989,-44952,-44915,
    -44879,-44842,-44806,-44769,-44732,-44695,-44659,-44622,
    -44585,-44548,-44511,-44474,-44437,-44400,-44363,-44326,
    -44289,-44252,-44215,-44178,-44141,-44104,-44067,-44029,
    -43992,-43955,-43918,-43880,-43843,-43806,-43768,-43731,
    -43693,-43656,-43618,-43581,-43543,-43506,-43468,-43430,
    -43393,-43355,-43317,-43280,-43242,-43204,-43166,-43128,
    -43091,-43053,-43015,-42977,-42939,-42901,-42863,-42825,
    -42787,-42749,-42711,-42672,-42634,-42596,-42558,-42520,
    -42481,-42443,-42405,-42366,-42328,-42290,-42251,-42213,
    -42174,-42136,-42097,-42059,-42020,-41982,-41943,-41904,
    -41866,-41827,-41788,-41750,-41711,-41672,-41633,-41595,
    -41556,-41517,-41478,-41439,-41400,-41361,-41322,-41283,
    -41244,-41205,-41166,-41127,-41087,-41048,-41009,-40970,
    -40931,-40891,-40852,-40813,-40773,-40734,-40695,-40655,
    -40616,-40576,-40537,-40497,-40458,-40418,-40379,-40339,
    -40299,-40260,-40220,-40180,-40141,-40101,-40061,-40021,
    -39982,-39942,-39902,-39862,-39822,-39782,-39742,-39702,
    -39662,-39622,-39582,-39542,-39502,-39462,-39422,-39382,
    -39341,-39301,-39261,-39221,-39180,-39140,-39100,-39059,
    -39019,-38979,-38938,-38898,-38857,-38817,-38776,-38736,
    -38695,-38655,-38614,-38573,-38533,-38492,-38451,-38411,
    -38370,-38329,-38288,-38248,-38207,-38166,-38125,-38084,
    -38043,-38002,-37961,-37920,-37879,-37838,-37797,-37756,
    -37715,-37674,-37633,-37592,-37550,-37509,-37468,-37427,
    -37386,-37344,-37303,-37262,-37220,-37179,-37137,-37096,
    -37055,-37013,-36972,-36930,-36889,-36847,-36805,-36764,
    -36722,-36681,-36639,-36597,-36556,-36514,-36472,-36430,
    -36388,-36347,-36305,-36263,-36221,-36179,-36137,-36095,
    -36053,-36011,-35969,-35927,-35885,-35843,-35801,-35759,
    -35717,-35675,-35633,-35590,-35548,-35506,-35464,-35421,
    -35379,-35337,-35294,-35252,-35210,-35167,-35125,-35082,
    -35040,-34997,-34955,-34912,-34870,-34827,-34785,-34742,
    -34699,-34657,-34614,-34571,-34529,-34486,-34443,-34400,
    -34358,-34315,-34272,-34229,-34186,-34143,-34100,-34057,
    -34015,-33972,-33929,-33886,-33843,-33799,-33756,-33713,
    -33670,-33627,-33584,-33541,-33498,-33454,-33411,-33368,
    -33325,-33281,-33238,-33195,-33151,-33108,-33065,-33021,
    -32978,-32934,-32891,-32847,-32804,-32760,-32717,-32673,
    -32630,-32586,-32542,-32499,-32455,-32411,-32368,-32324,
    -32280,-32236,-32193,-32149,-32105,-32061,-32017,-31974,
    -31930,-31886,-31842,-31798,-31754,-31710,-31666,-31622,
    -31578,-31534,-31490,-31446,-31402,-31357,-31313,-31269,
    -31225,-31181,-31136,-31092,-31048,-31004,-30959,-30915,
    -30871,-30826,-30782,-30738,-30693,-30649,-30604,-30560,
    -30515,-30471,-30426,-30382,-30337,-30293,-30248,-30204,
    -30159,-30114,-30070,-30025,-29980,-29936,-29891,-29846,
    -29801,-29757,-29712,-29667,-29622,-29577,-29533,-29488,
    -29443,-29398,-29353,-29308,-29263,-29218,-29173,-29128,
    -29083,-29038,-28993,-28948,-28903,-28858,-28812,-28767,
    -28722,-28677,-28632,-28586,-28541,-28496,-28451,-28405,
    -28360,-28315,-28269,-28224,-28179,-28133,-28088,-28042,
    -27997,-27952,-27906,-27861,-27815,-27770,-27724,-27678,
    -27633,-27587,-27542,-27496,-27450,-27405,-27359,-27313,
    -27268,-27222,-27176,-27131,-27085,-27039,-26993,-26947,
    -26902,-26856,-26810,-26764,-26718,-26672,-26626,-26580,
    -26534,-26488,-26442,-26396,-26350,-26304,-26258,-26212,
    -26166,-26120,-26074,-26028,-25982,-25936,-25889,-25843,
    -25797,-25751,-25705,-25658,-25612,-25566,-25520,-25473,
    -25427,-25381,-25334,-25288,-25241,-25195,-25149,-25102,
    -25056,-25009,-24963,-24916,-24870,-24823,-24777,-24730,
    -24684,-24637,-24591,-24544,-24497,-24451,-24404,-24357,
    -24311,-24264,-24217,-24171,-24124,-24077,-24030,-23984,
    -23937,-23890,-23843,-23796,-23750,-23703,-23656,-23609,
    -23562,-23515,-23468,-23421,-23374,-23327,-23280,-23233,
    -23186,-23139,-23092,-23045,-22998,-22951,-22904,-22857,
    -22810,-22763,-22716,-22668,-22621,-22574,-22527,-22480,
    -22432,-22385,-22338,-22291,-22243,-22196,-22149,-22102,
    -22054,-22007,-21960,-21912,-21865,-21817,-21770,-21723,
    -21675,-21628,-21580,-21533,-21485,-21438,-21390,-21343,
    -21295,-21248,-21200,-21153,-21105,-21057,-21010,-20962,
    -20915,-20867,-20819,-20772,-20724,-20676,-20629,-20581,
    -20533,-20485,-20438,-20390,-20342,-20294,-20246,-20199,
    -20151,-20103,-20055,-20007,-19959,-19912,-19864,-19816,
    -19768,-19720,-19672,-19624,-19576,-19528,-19480,-19432,
    -19384,-19336,-19288,-19240,-19192,-19144,-19096,-19048,
    -19000,-18951,-18903,-18855,-18807,-18759,-18711,-18663,
    -18614,-18566,-18518,-18470,-18421,-18373,-18325,-18277,
    -18228,-18180,-18132,-18084,-18035,-17987,-17939,-17890,
    -17842,-17793,-17745,-17697,-17648,-17600,-17551,-17503,
    -17455,-17406,-17358,-17309,-17261,-17212,-17164,-17115,
    -17067,-17018,-16970,-16921,-16872,-16824,-16775,-16727,
    -16678,-16629,-16581,-16532,-16484,-16435,-16386,-16338,
    -16289,-16240,-16191,-16143,-16094,-16045,-15997,-15948,
    -15899,-15850,-15802,-15753,-15704,-15655,-15606,-15557,
    -15509,-15460,-15411,-15362,-15313,-15264,-15215,-15167,
    -15118,-15069,-15020,-14971,-14922,-14873,-14824,-14775,
    -14726,-14677,-14628,-14579,-14530,-14481,-14432,-14383,
    -14334,-14285,-14236,-14187,-14138,-14089,-14040,-13990,
    -13941,-13892,-13843,-13794,-13745,-13696,-13647,-13597,
    -13548,-13499,-13450,-13401,-13351,-13302,-13253,-13204,
    -13154,-13105,-13056,-13007,-12957,-12908,-12859,-12810,
    -12760,-12711,-12662,-12612,-12563,-12514,-12464,-12415,
    -12366,-12316,-12267,-12217,-12168,-12119,-12069,-12020,
    -11970,-11921,-11872,-11822,-11773,-11723,-11674,-11624,
    -11575,-11525,-11476,-11426,-11377,-11327,-11278,-11228,
    -11179,-11129,-11080,-11030,-10981,-10931,-10882,-10832,
    -10782,-10733,-10683,-10634,-10584,-10534,-10485,-10435,
    -10386,-10336,-10286,-10237,-10187,-10137,-10088,-10038,
    -9988,-9939,-9889,-9839,-9790,-9740,-9690,-9640,
    -9591,-9541,-9491,-9442,-9392,-9342,-9292,-9243,
    -9193,-9143,-9093,-9043,-8994,-8944,-8894,-8844,
    -8794,-8745,-8695,-8645,-8595,-8545,-8496,-8446,
    -8396,-8346,-8296,-8246,-8196,-8147,-8097,-8047,
    -7997,-7947,-7897,-7847,-7797,-7747,-7697,-7648,
    -7598,-7548,-7498,-7448,-7398,-7348,-7298,-7248,
    -7198,-7148,-7098,-7048,-6998,-6948,-6898,-6848,
    -6798,-6748,-6698,-6648,-6598,-6548,-6498,-6448,
    -6398,-6348,-6298,-6248,-6198,-6148,-6098,-6048,
    -5998,-5948,-5898,-5848,-5798,-5747,-5697,-5647,
    -5597,-5547,-5497,-5447,-5397,-5347,-5297,-5247,
    -5197,-5146,-5096,-5046,-4996,-4946,-4896,-4846,
    -4796,-4745,-4695,-4645,-4595,-4545,-4495,-4445,
    -4394,-4344,-4294,-4244,-4194,-4144,-4093,-4043,
    -3993,-3943,-3893,-3843,-3792,-3742,-3692,-3642,
    -3592,-3541,-3491,-3441,-3391,-3341,-3291,-3240,
    -3190,-3140,-3090,-3039,-2989,-2939,-2889,-2839,
    -2788,-2738,-2688,-2638,-2588,-2537,-2487,-2437,
    -2387,-2336,-2286,-2236,-2186,-2135,-2085,-2035,
    -1985,-1934,-1884,-1834,-1784,-1733,-1683,-1633,
    -1583,-1532,-1482,-1432,-1382,-1331,-1281,-1231,
    -1181,-1130,-1080,-1030,-980,-929,-879,-829,
    -779,-728,-678,-628,-578,-527,-477,-427,
    -376,-326,-276,-226,-175,-125,-75,-25,
    25,75,125,175,226,276,326,376,
    427,477,527,578,628,678,728,779,
    829,879,929,980,1030,1080,1130,1181,
    1231,1281,1331,1382,1432,1482,1532,1583,
    1633,1683,1733,1784,1834,1884,1934,1985,
    2035,2085,2135,2186,2236,2286,2336,2387,
    2437,2487,2537,2587,2638,2688,2738,2788,
    2839,2889,2939,2989,3039,3090,3140,3190,
    3240,3291,3341,3391,3441,3491,3542,3592,
    3642,3692,3742,3792,3843,3893,3943,3993,
    4043,4093,4144,4194,4244,4294,4344,4394,
    4445,4495,4545,4595,4645,4695,4745,4796,
    4846,4896,4946,4996,5046,5096,5146,5197,
    5247,5297,5347,5397,5447,5497,5547,5597,
    5647,5697,5747,5798,5848,5898,5948,5998,
    6048,6098,6148,6198,6248,6298,6348,6398,
    6448,6498,6548,6598,6648,6698,6748,6798,
    6848,6898,6948,6998,7048,7098,7148,7198,
    7248,7298,7348,7398,7448,7498,7548,7598,
    7648,7697,7747,7797,7847,7897,7947,7997,
    8047,8097,8147,8196,8246,8296,8346,8396,
    8446,8496,8545,8595,8645,8695,8745,8794,
    8844,8894,8944,8994,9043,9093,9143,9193,
    9243,9292,9342,9392,9442,9491,9541,9591,
    9640,9690,9740,9790,9839,9889,9939,9988,
    10038,10088,10137,10187,10237,10286,10336,10386,
    10435,10485,10534,10584,10634,10683,10733,10782,
    10832,10882,10931,10981,11030,11080,11129,11179,
    11228,11278,11327,11377,11426,11476,11525,11575,
    11624,11674,11723,11773,11822,11872,11921,11970,
    12020,12069,12119,12168,12218,12267,12316,12366,
    12415,12464,12514,12563,12612,12662,12711,12760,
    12810,12859,12908,12957,13007,13056,13105,13154,
    13204,13253,13302,13351,13401,13450,13499,13548,
    13597,13647,13696,13745,13794,13843,13892,13941,
    13990,14040,14089,14138,14187,14236,14285,14334,
    14383,14432,14481,14530,14579,14628,14677,14726,
    14775,14824,14873,14922,14971,15020,15069,15118,
    15167,15215,15264,15313,15362,15411,15460,15509,
    15557,15606,15655,15704,15753,15802,15850,15899,
    15948,15997,16045,16094,16143,16191,16240,16289,
    16338,16386,16435,16484,16532,16581,16629,16678,
    16727,16775,16824,16872,16921,16970,17018,17067,
    17115,17164,17212,17261,17309,17358,17406,17455,
    17503,17551,17600,17648,17697,17745,17793,17842,
    17890,17939,17987,18035,18084,18132,18180,18228,
    18277,18325,18373,18421,18470,18518,18566,18614,
    18663,18711,18759,18807,18855,18903,18951,19000,
    19048,19096,19144,19192,19240,19288,19336,19384,
    19432,19480,19528,19576,19624,19672,19720,19768,
    19816,19864,19912,19959,20007,20055,20103,20151,
    20199,20246,20294,20342,20390,20438,20485,20533,
    20581,20629,20676,20724,20772,20819,20867,20915,
    20962,21010,21057,21105,21153,21200,21248,21295,
    21343,21390,21438,21485,21533,21580,21628,21675,
    21723,21770,21817,21865,21912,21960,22007,22054,
    22102,22149,22196,22243,22291,22338,22385,22432,
    22480,22527,22574,22621,22668,22716,22763,22810,
    22857,22904,22951,22998,23045,23092,23139,23186,
    23233,23280,23327,23374,23421,23468,23515,23562,
    23609,23656,23703,23750,23796,23843,23890,23937,
    23984,24030,24077,24124,24171,24217,24264,24311,
    24357,24404,24451,24497,24544,24591,24637,24684,
    24730,24777,24823,24870,24916,24963,25009,25056,
    25102,25149,25195,25241,25288,25334,25381,25427,
    25473,25520,25566,25612,25658,25705,25751,25797,
    25843,25889,25936,25982,26028,26074,26120,26166,
    26212,26258,26304,26350,26396,26442,26488,26534,
    26580,26626,26672,26718,26764,26810,26856,26902,
    26947,26993,27039,27085,27131,27176,27222,27268,
    27313,27359,27405,27450,27496,27542,27587,27633,
    27678,27724,27770,27815,27861,27906,27952,27997,
    28042,28088,28133,28179,28224,28269,28315,28360,
    28405,28451,28496,28541,28586,28632,28677,28722,
    28767,28812,28858,28903,28948,28993,29038,29083,
    29128,29173,29218,29263,29308,29353,29398,29443,
    29488,29533,29577,29622,29667,29712,29757,29801,
    29846,29891,29936,29980,30025,30070,30114,30159,
    30204,30248,30293,30337,30382,30427,30471,30516,
    30560,30604,30649,30693,30738,30782,30826,30871,
    30915,30959,31004,31048,31092,31136,31181,31225,
    31269,31313,31357,31402,31446,31490,31534,31578,
    31622,31666,31710,31754,31798,31842,31886,31930,
    31974,32017,32061,32105,32149,32193,32236,32280,
    32324,32368,32411,32455,32499,32542,32586,32630,
    32673,32717,32760,32804,32847,32891,32934,32978,
    33021,33065,33108,33151,33195,33238,33281,33325,
    33368,33411,33454,33498,33541,33584,33627,33670,
    33713,33756,33799,33843,33886,33929,33972,34015,
    34057,34100,34143,34186,34229,34272,34315,34358,
    34400,34443,34486,34529,34571,34614,34657,34699,
    34742,34785,34827,34870,34912,34955,34997,35040,
    35082,35125,35167,35210,35252,35294,35337,35379,
    35421,35464,35506,35548,35590,35633,35675,35717,
    35759,35801,35843,35885,35927,35969,36011,36053,
    36095,36137,36179,36221,36263,36305,36347,36388,
    36430,36472,36514,36556,36597,36639,36681,36722,
    36764,36805,36847,36889,36930,36972,37013,37055,
    37096,37137,37179,37220,37262,37303,37344,37386,
    37427,37468,37509,37551,37592,37633,37674,37715,
    37756,37797,37838,37879,37920,37961,38002,38043,
    38084,38125,38166,38207,38248,38288,38329,38370,
    38411,38451,38492,38533,38573,38614,38655,38695,
    38736,38776,38817,38857,38898,38938,38979,39019,
    39059,39100,39140,39180,39221,39261,39301,39341,
    39382,39422,39462,39502,39542,39582,39622,39662,
    39702,39742,39782,39822,39862,39902,39942,39982,
    40021,40061,40101,40141,40180,40220,40260,40299,
    40339,40379,40418,40458,40497,40537,40576,40616,
    40655,40695,40734,40773,40813,40852,40891,40931,
    40970,41009,41048,41087,41127,41166,41205,41244,
    41283,41322,41361,41400,41439,41478,41517,41556,
    41595,41633,41672,41711,41750,41788,41827,41866,
    41904,41943,41982,42020,42059,42097,42136,42174,
    42213,42251,42290,42328,42366,42405,42443,42481,
    42520,42558,42596,42634,42672,42711,42749,42787,
    42825,42863,42901,42939,42977,43015,43053,43091,
    43128,43166,43204,43242,43280,43317,43355,43393,
    43430,43468,43506,43543,43581,43618,43656,43693,
    43731,43768,43806,43843,43880,43918,43955,43992,
    44029,44067,44104,44141,44178,44215,44252,44289,
    44326,44363,44400,44437,44474,44511,44548,44585,
    44622,44659,44695,44732,44769,44806,44842,44879,
    44915,44952,44989,45025,45062,45098,45135,45171,
    45207,45244,45280,45316,45353,45389,45425,45462,
    45498,45534,45570,45606,45642,45678,45714,45750,
    45786,45822,45858,45894,45930,45966,46002,46037,
    46073,46109,46145,46180,46216,46252,46287,46323,
    46358,46394,46429,46465,46500,46536,46571,46606,
    46642,46677,46712,46747,46783,46818,46853,46888,
    46923,46958,46993,47028,47063,47098,47133,47168,
    47203,47238,47273,47308,47342,47377,47412,47446,
    47481,47516,47550,47585,47619,47654,47688,47723,
    47757,47792,47826,47861,47895,47929,47963,47998,
    48032,48066,48100,48134,48168,48202,48237,48271,
    48305,48338,48372,48406,48440,48474,48508,48542,
    48575,48609,48643,48676,48710,48744,48777,48811,
    48844,48878,48911,48945,48978,49012,49045,49078,
    49112,49145,49178,49211,49244,49278,49311,49344,
    49377,49410,49443,49476,49509,49542,49575,49608,
    49640,49673,49706,49739,49771,49804,49837,49869,
    49902,49935,49967,50000,50032,50064,50097,50129,
    50162,50194,50226,50259,50291,50323,50355,50387,
    50420,50452,50484,50516,50548,50580,50612,50644,
    50675,50707,50739,50771,50803,50834,50866,50898,
    50929,50961,50993,51024,51056,51087,51119,51150,
    51182,51213,51244,51276,51307,51338,51369,51401,
    51432,51463,51494,51525,51556,51587,51618,51649,
    51680,51711,51742,51773,51803,51834,51865,51896,
    51926,51957,51988,52018,52049,52079,52110,52140,
    52171,52201,52231,52262,52292,52322,52353,52383,
    52413,52443,52473,52503,52534,52564,52594,52624,
    52653,52683,52713,52743,52773,52803,52832,52862,
    52892,52922,52951,52981,53010,53040,53069,53099,
    53128,53158,53187,53216,53246,53275,53304,53334,
    53363,53392,53421,53450,53479,53508,53537,53566,
    53595,53624,53653,53682,53711,53739,53768,53797,
    53826,53854,53883,53912,53940,53969,53997,54026,
    54054,54082,54111,54139,54167,54196,54224,54252,
    54280,54309,54337,54365,54393,54421,54449,54477,
    54505,54533,54560,54588,54616,54644,54672,54699,
    54727,54755,54782,54810,54837,54865,54892,54920,
    54947,54974,55002,55029,55056,55084,55111,55138,
    55165,55192,55219,55246,55274,55300,55327,55354,
    55381,55408,55435,55462,55489,55515,55542,55569,
    55595,55622,55648,55675,55701,55728,55754,55781,
    55807,55833,55860,55886,55912,55938,55965,55991,
    56017,56043,56069,56095,56121,56147,56173,56199,
    56225,56250,56276,56302,56328,56353,56379,56404,
    56430,56456,56481,56507,56532,56557,56583,56608,
    56633,56659,56684,56709,56734,56760,56785,56810,
    56835,56860,56885,56910,56935,56959,56984,57009,
    57034,57059,57083,57108,57133,57157,57182,57206,
    57231,57255,57280,57304,57329,57353,57377,57402,
    57426,57450,57474,57498,57522,57546,57570,57594,
    57618,57642,57666,57690,57714,57738,57762,57785,
    57809,57833,57856,57880,57903,57927,57950,57974,
    57997,58021,58044,58067,58091,58114,58137,58160,
    58183,58207,58230,58253,58276,58299,58322,58345,
    58367,58390,58413,58436,58459,58481,58504,58527,
    58549,58572,58594,58617,58639,58662,58684,58706,
    58729,58751,58773,58795,58818,58840,58862,58884,
    58906,58928,58950,58972,58994,59016,59038,59059,
    59081,59103,59125,59146,59168,59190,59211,59233,
    59254,59276,59297,59318,59340,59361,59382,59404,
    59425,59446,59467,59488,59509,59530,59551,59572,
    59593,59614,59635,59656,59677,59697,59718,59739,
    59759,59780,59801,59821,59842,59862,59883,59903,
    59923,59944,59964,59984,60004,60025,60045,60065,
    60085,60105,60125,60145,60165,60185,60205,60225,
    60244,60264,60284,60304,60323,60343,60363,60382,
    60402,60421,60441,60460,60479,60499,60518,60537,
    60556,60576,60595,60614,60633,60652,60671,60690,
    60709,60728,60747,60766,60785,60803,60822,60841,
    60859,60878,60897,60915,60934,60952,60971,60989,
    61007,61026,61044,61062,61081,61099,61117,61135,
    61153,61171,61189,61207,61225,61243,61261,61279,
    61297,61314,61332,61350,61367,61385,61403,61420,
    61438,61455,61473,61490,61507,61525,61542,61559,
    61577,61594,61611,61628,61645,61662,61679,61696,
    61713,61730,61747,61764,61780,61797,61814,61831,
    61847,61864,61880,61897,61913,61930,61946,61963,
    61979,61995,62012,62028,62044,62060,62076,62092,
    62108,62125,62141,62156,62172,62188,62204,62220,
    62236,62251,62267,62283,62298,62314,62329,62345,
    62360,62376,62391,62407,62422,62437,62453,62468,
    62483,62498,62513,62528,62543,62558,62573,62588,
    62603,62618,62633,62648,62662,62677,62692,62706,
    62721,62735,62750,62764,62779,62793,62808,62822,
    62836,62850,62865,62879,62893,62907,62921,62935,
    62949,62963,62977,62991,63005,63019,63032,63046,
    63060,63074,63087,63101,63114,63128,63141,63155,
    63168,63182,63195,63208,63221,63235,63248,63261,
    63274,63287,63300,63313,63326,63339,63352,63365,
    63378,63390,63403,63416,63429,63441,63454,63466,
    63479,63491,63504,63516,63528,63541,63553,63565,
    63578,63590,63602,63614,63626,63638,63650,63662,
    63674,63686,63698,63709,63721,63733,63745,63756,
    63768,63779,63791,63803,63814,63825,63837,63848,
    63859,63871,63882,63893,63904,63915,63927,63938,
    63949,63960,63971,63981,63992,64003,64014,64025,
    64035,64046,64057,64067,64078,64088,64099,64109,
    64120,64130,64140,64151,64161,64171,64181,64192,
    64202,64212,64222,64232,64242,64252,64261,64271,
    64281,64291,64301,64310,64320,64330,64339,64349,
    64358,64368,64377,64387,64396,64405,64414,64424,
    64433,64442,64451,64460,64469,64478,64487,64496,
    64505,64514,64523,64532,64540,64549,64558,64566,
    64575,64584,64592,64600,64609,64617,64626,64634,
    64642,64651,64659,64667,64675,64683,64691,64699,
    64707,64715,64723,64731,64739,64747,64754,64762,
    64770,64777,64785,64793,64800,64808,64815,64822,
    64830,64837,64844,64852,64859,64866,64873,64880,
    64887,64895,64902,64908,64915,64922,64929,64936,
    64943,64949,64956,64963,64969,64976,64982,64989,
    64995,65002,65008,65015,65021,65027,65033,65040,
    65046,65052,65058,65064,65070,65076,65082,65088,
    65094,65099,65105,65111,65117,65122,65128,65133,
    65139,65144,65150,65155,65161,65166,65171,65177,
    65182,65187,65192,65197,65202,65207,65212,65217,
    65222,65227,65232,65237,65242,65246,65251,65256,
    65260,65265,65270,65274,65279,65283,65287,65292,
    65296,65300,65305,65309,65313,65317,65321,65325,
    65329,65333,65337,65341,65345,65349,65352,65356,
    65360,65363,65367,65371,65374,65378,65381,65385,
    65388,65391,65395,65398,65401,65404,65408,65411,
    65414,65417,65420,65423,65426,65429,65431,65434,
    65437,65440,65442,65445,65448,65450,65453,65455,
    65458,65460,65463,65465,65467,65470,65472,65474,
    65476,65478,65480,65482,65484,65486,65488,65490,
    65492,65494,65496,65497,65499,65501,65502,65504,
    65505,65507,65508,65510,65511,65513,65514,65515,
    65516,65518,65519,65520,65521,65522,65523,65524,
    65525,65526,65527,65527,65528,65529,65530,65530,
    65531,65531,65532,65532,65533,65533,65534,65534,
    65534,65535,65535,65535,65535,65535,65535,65535
)]!

const finecosine = unsafe { &finesine[fineangles / 4] }

const fineangles = 10240
