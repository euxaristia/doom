@[translated]
module main

// Network struct read/write support: placeholder manual port.
