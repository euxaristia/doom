module core

pub fn r_draw() {}
