module core

pub fn deh_frame_init() {}
