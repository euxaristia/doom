@[translated]
module main

// OPL3 core: placeholder manual port.
