@[translated]
module main

// Setup icon data: placeholder manual port.
