@[has_globals]
module core

__global deh_frame_overrides = 0

pub fn deh_frame_init() {
	deh_frame_overrides = 0
}
