@[translated]
module main

// OPL droplay example: placeholder manual port.
