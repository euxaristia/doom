@[translated]
module main

// Dedicated networking support: placeholder manual port.
