@[translated]
module main

// Textscreen file select widget: placeholder manual port.
