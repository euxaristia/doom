module core

pub fn p_doors_do_door_stub(line &Line, doortype int) int {
	_ = line
	_ = doortype
	return 0
}

pub fn p_doors_vertical_door_stub(line &Line, mobj &Mobj) {
	_ = line
	_ = mobj
}
