@[translated]
module main

// Disk icon module: placeholder manual port.
