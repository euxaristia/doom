module core

// Networking stubs; full netcode is not wired yet.
pub fn d_net_init() {}
pub fn d_net_shutdown() {}
pub fn d_net_connect() bool { return false }
pub fn d_net_disconnect() {}
