@[translated]
module main

// Setup mode module: placeholder manual port.
