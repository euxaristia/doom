module core

pub fn r_init() {}
