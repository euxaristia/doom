@[translated]
module main

// High-resolution video hooks: placeholder manual port.
