@[translated]
module main

// Video primitives module: placeholder manual port.
