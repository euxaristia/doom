module core

pub fn deh_weapon_init() {}
