@[has_globals]
module core

__global deh_sound_overrides = 0

pub fn deh_sound_init() {
	deh_sound_overrides = 0
}
