@[translated]
module main

// Textscreen spin control widget: placeholder manual port.
