@[translated]
module main

// Setup sound module: placeholder manual port.
