module core

pub fn p_check_sight_stub(t1 &Mobj, t2 &Mobj) bool {
	_ = t1
	_ = t2
	return true
}
