@[translated]
module main

// Network packet support: placeholder manual port.
