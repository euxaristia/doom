@[translated]
module main

// Digital music pack support: placeholder manual port.
