@[translated]
module main

// Setup main menu module: placeholder manual port.
