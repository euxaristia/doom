@[translated]
module main

// OPL music support: placeholder manual port.
