@[translated]
module main

// Window icon data is omitted in this minimal manual port.
