@[translated]
module main

// Textscreen strut widget: placeholder manual port.
