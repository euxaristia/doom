module core

// Carries out all thinking of monsters and players.
pub fn p_ticker() {}
