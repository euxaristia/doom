module main

@[weak] __global ( test_array [3]int )

fn main() {
    // This is just a test
}