module core

pub fn p_ceilng_do_ceiling_stub(line &Line, ceilingtype int) int {
	_ = line
	_ = ceilingtype
	return 0
}
