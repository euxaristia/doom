@[has_globals]
module core

__global deh_cheats_applied = false

pub fn deh_cheat_init() {
	deh_cheats_applied = false
}
