@[translated]
module main

// Setup textscreen joystick axis module: placeholder manual port.
