@[translated]
module main

// OPL SDL backend: placeholder manual port.
