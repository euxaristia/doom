@[translated]
module main

// Textscreen dropdown widget: placeholder manual port.
