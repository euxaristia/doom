module core

pub fn p_give_power(player voidptr, power int) bool {
	_ = player
	_ = power
	return false
}
