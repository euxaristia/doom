module core

pub fn p_move_player(player &Player) {
	_ = player
}

pub fn p_calc_height(player &Player) {
	_ = player
}
