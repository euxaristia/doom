@[translated]
module main

// Textscreen GUI core: placeholder manual port.
