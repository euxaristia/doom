module core

pub fn p_lights_turn_on_stub(line &Line, bright int) {
	_ = line
	_ = bright
}

pub fn p_lights_start_strobing_stub(line &Line) {
	_ = line
}
