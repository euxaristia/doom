@[translated]
module main

// Textscreen separator widget: placeholder manual port.
