@[translated]
module main

// Setup mouse module: placeholder manual port.
