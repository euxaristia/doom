module core

pub fn p_approx_distance(dx Fixed, dy Fixed) Fixed {
	_ = dx
	_ = dy
	return 0
}
