module core

// Minimal renderer data placeholders.
pub fn r_init_data() {}
