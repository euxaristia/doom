@[translated]
module main

// Network I/O support: placeholder manual port.
