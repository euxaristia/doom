@[translated]
module main

// Network GUI support: placeholder manual port.
