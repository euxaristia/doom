@[has_globals]
module core

__global deh_weapon_overrides = 0

pub fn deh_weapon_init() {
	deh_weapon_overrides = 0
}
