@[translated]
module main

// OPL OpenBSD backend: placeholder manual port.
