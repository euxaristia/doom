module core

pub struct CheatSeq {
pub mut:
	sequence string
}
