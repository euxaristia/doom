@[translated]
module main

// Setup keyboard module: placeholder manual port.
