@[translated]
module main

// Textscreen calculator example: placeholder manual port.
