@[translated]
module main

// SDL music backend: placeholder manual port.
