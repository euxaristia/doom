module core

pub struct Mobj {
pub mut:
	thinker Thinker
}
