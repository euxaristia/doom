@[translated]
module main

// OPL ioperm syscalls: placeholder manual port.
