module core

// Minimal English string placeholders.
pub const presskey = 'press a key'
