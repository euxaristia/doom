@[translated]
module main

// OPL timer: placeholder manual port.
