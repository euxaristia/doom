module core

pub fn r_render_bsp() {}
