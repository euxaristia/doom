@[translated]
module main

// Textscreen UTF-8 helpers: placeholder manual port.
