@[translated]
module main

// Network petname support: placeholder manual port.
