@[translated]
module main

// stdio WAD file backend: placeholder manual port.
