@[translated]
module main

// Setup display module: placeholder manual port.
