@[translated]
module main

// Setup compatibility module: placeholder manual port.
