@[translated]
module main

// MIDI file parsing: placeholder manual port.
