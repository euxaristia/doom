@[translated]
module main

// Setup execute module: placeholder manual port.
