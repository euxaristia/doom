@[translated]
module main

// MIDI pipe support: placeholder manual port.
