@[translated]
module main

// Textscreen button widget: placeholder manual port.
