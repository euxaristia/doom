@[has_globals]
module core

__global deh_thing_overrides = 0

pub fn deh_thing_init() {
	deh_thing_overrides = 0
}
