@[translated]
module main

// Joystick binding and init hooks.

@[export: 'I_BindJoystickVariables']
pub fn i_bind_joystick_variables() {
	// No-op placeholder.
}

@[export: 'I_InitJoystick']
pub fn i_init_joystick() {
	// No-op placeholder.
}
