@[translated]
module main

// OPL Linux backend: placeholder manual port.
