module core

pub struct NetConnectData {}

pub struct NetGameSettings {}
