@[translated]
module main

// OPL Win32 backend: placeholder manual port.
